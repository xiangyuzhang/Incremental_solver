
module c2670 (N1,N2,N3,N4,N5,N6,N7,N8,N11,N14,
              N15,N16,N19,N20,N21,N22,N23,N24,N25,N26,
              N27,N28,N29,N32,N33,N34,N35,N36,N37,N40,
              N43,N44,N47,N48,N49,N50,N51,N52,N53,N54,
              N55,N56,N57,N60,N61,N62,N63,N64,N65,N66,
              N67,N68,N69,N72,N73,N74,N75,N76,N77,N78,
              N79,N80,N81,N82,N85,N86,N87,N88,N89,N90,
              N91,N92,N93,N94,N95,N96,N99,N100,N101,N102,
              N103,N104,N105,N106,N107,N108,N111,N112,N113,N114,
              N115,N116,N117,N118,N119,N120,N123,N124,N125,N126,
              N127,N128,N129,N130,N131,N132,N135,N136,N137,N138,
              N139,N140,N141,N142,N219,N224,N227,N230,N231,N234,
              N237,N241,N246,N253,N256,N259,N262,N263,N266,N269,
              N272,N275,N278,N281,N284,N287,N290,N294,N297,N301,
              N305,N309,N313,N316,N319,N322,N325,N328,N331,N334,
              N337,N340,N343,N346,N349,N352,N355,N143_I,N144_I,N145_I,
              N146_I,N147_I,N148_I,N149_I,N150_I,N151_I,N152_I,N153_I,N154_I,N155_I,
              N156_I,N157_I,N158_I,N159_I,N160_I,N161_I,N162_I,N163_I,N164_I,N165_I,
              N166_I,N167_I,N168_I,N169_I,N170_I,N171_I,N172_I,N173_I,N174_I,N175_I,
              N176_I,N177_I,N178_I,N179_I,N180_I,N181_I,N182_I,N183_I,N184_I,N185_I,
              N186_I,N187_I,N188_I,N189_I,N190_I,N191_I,N192_I,N193_I,N194_I,N195_I,
              N196_I,N197_I,N198_I,N199_I,N200_I,N201_I,N202_I,N203_I,N204_I,N205_I,
              N206_I,N207_I,N208_I,N209_I,N210_I,N211_I,N212_I,N213_I,N214_I,N215_I,
              N216_I,N217_I,N218_I,N398,N400,N401,N419,N420,N456,N457,
              N458,N487,N488,N489,N490,N491,N492,N493,N494,N792,
              N799,N805,N1026,N1028,N1029,N1269,N1277,N1448,N1726,N1816,
              N1817,N1818,N1819,N1820,N1821,N1969,N1970,N1971,N2010,N2012,
              N2014,N2016,N2018,N2020,N2022,N2387,N2388,N2389,N2390,N2496,
              N2643,N2644,N2891,N2925,N2970,N2971,N3038,N3079,N3546,N3671,
              N3803,N3804,N3809,N3851,N3875,N3881,N3882,N143_O,N144_O,N145_O,
              N146_O,N147_O,N148_O,N149_O,N150_O,N151_O,N152_O,N153_O,N154_O,N155_O,
              N156_O,N157_O,N158_O,N159_O,N160_O,N161_O,N162_O,N163_O,N164_O,N165_O,
              N166_O,N167_O,N168_O,N169_O,N170_O,N171_O,N172_O,N173_O,N174_O,N175_O,
              N176_O,N177_O,N178_O,N179_O,N180_O,N181_O,N182_O,N183_O,N184_O,N185_O,
              N186_O,N187_O,N188_O,N189_O,N190_O,N191_O,N192_O,N193_O,N194_O,N195_O,
              N196_O,N197_O,N198_O,N199_O,N200_O,N201_O,N202_O,N203_O,N204_O,N205_O,
              N206_O,N207_O,N208_O,N209_O,N210_O,N211_O,N212_O,N213_O,N214_O,N215_O,
              N216_O,N217_O,N218_O);

input N1,N2,N3,N4,N5,N6,N7,N8,N11,N14,
      N15,N16,N19,N20,N21,N22,N23,N24,N25,N26,
      N27,N28,N29,N32,N33,N34,N35,N36,N37,N40,
      N43,N44,N47,N48,N49,N50,N51,N52,N53,N54,
      N55,N56,N57,N60,N61,N62,N63,N64,N65,N66,
      N67,N68,N69,N72,N73,N74,N75,N76,N77,N78,
      N79,N80,N81,N82,N85,N86,N87,N88,N89,N90,
      N91,N92,N93,N94,N95,N96,N99,N100,N101,N102,
      N103,N104,N105,N106,N107,N108,N111,N112,N113,N114,
      N115,N116,N117,N118,N119,N120,N123,N124,N125,N126,
      N127,N128,N129,N130,N131,N132,N135,N136,N137,N138,
      N139,N140,N141,N142,N219,N224,N227,N230,N231,N234,
      N237,N241,N246,N253,N256,N259,N262,N263,N266,N269,
      N272,N275,N278,N281,N284,N287,N290,N294,N297,N301,
      N305,N309,N313,N316,N319,N322,N325,N328,N331,N334,
      N337,N340,N343,N346,N349,N352,N355,N143_I,N144_I,N145_I,
      N146_I,N147_I,N148_I,N149_I,N150_I,N151_I,N152_I,N153_I,N154_I,N155_I,
      N156_I,N157_I,N158_I,N159_I,N160_I,N161_I,N162_I,N163_I,N164_I,N165_I,
      N166_I,N167_I,N168_I,N169_I,N170_I,N171_I,N172_I,N173_I,N174_I,N175_I,
      N176_I,N177_I,N178_I,N179_I,N180_I,N181_I,N182_I,N183_I,N184_I,N185_I,
      N186_I,N187_I,N188_I,N189_I,N190_I,N191_I,N192_I,N193_I,N194_I,N195_I,
      N196_I,N197_I,N198_I,N199_I,N200_I,N201_I,N202_I,N203_I,N204_I,N205_I,
      N206_I,N207_I,N208_I,N209_I,N210_I,N211_I,N212_I,N213_I,N214_I,N215_I,
      N216_I,N217_I,N218_I ;

input   p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,
        p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,
        p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,
        p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,
        p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,
        p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,
        p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,
        p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,
        p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,
        p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,
        p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,
        p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,
        p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,
        p131,p132,p133,p134,p135,p136,p137,p138,p139,p140,
        p141,p142,p143,p144,p145,p146,p147,p148,p149,p150,
        p151,p152,p153,p154,p155,p156,p157,p158,p159,p160,
        p161,p162,p163,p164,p165,p166,p167,p168,p169,p170,
        p171,p172,p173,p174,p175,p176,p177,p178,p179,p180,
        p181,p182,p183,p184,p185,p186,p187,p188,p189,p190,
        p191,p192,p193,p194,p195,p196,p197,p198,p199,p200,
        p201,p202,p203,p204,p205,p206,p207,p208,p209,p210,
        p211,p212,p213,p214,p215,p216,p217,p218,p219,p220,
        p221,p222,p223,p224,p225,p226,p227,p228,p229,p230,
        p231,p232,p233,p234,p235,p236,p237,p238,p239,p240,
        p241,p242,p243,p244,p245,p246,p247,p248,p249,p250,
        p251,p252,p253,p254,p255,p256,p257,p258,p259,p260,
        p261,p262,p263,p264,p265,p266,p267,p268,p269,p270,
        p271,p272,p273,p274,p275,p276,p277,p278,p279,p280,
        p281,p282,p283,p284,p285,p286,p287,p288,p289,p290,
        p291,p292,p293,p294,p295,p296,p297,p298,p299,p300,
        p301,p302,p303,p304,p305,p306,p307,p308,p309,p310,
        p311,p312,p313,p314,p315,p316,p317,p318,p319,p320,
        p321,p322,p323,p324,p325,p326,p327,p328,p329,p330,
        p331,p332,p333,p334,p335,p336,p337,p338,p339,p340,
        p341,p342,p343,p344,p345,p346,p347,p348,p349,p350,
        p351,p352,p353,p354,p355,p356,p357,p358,p359,p360,
        p361,p362,p363,p364,p365,p366,p367,p368,p369,p370,
        p371,p372,p373,p374,p375,p376,p377,p378,p379,p380 ;

output N398,N400,N401,N419,N420,N456,N457,N458,N487,N488,
       N489,N490,N491,N492,N493,N494,N792,N799,N805,N1026,
       N1028,N1029,N1269,N1277,N1448,N1726,N1816,N1817,N1818,N1819,
       N1820,N1821,N1969,N1970,N1971,N2010,N2012,N2014,N2016,N2018,
       N2020,N2022,N2387,N2388,N2389,N2390,N2496,N2643,N2644,N2891,
       N2925,N2970,N2971,N3038,N3079,N3546,N3671,N3803,N3804,N3809,
       N3851,N3875,N3881,N3882,N143_O,N144_O,N145_O,N146_O,N147_O,N148_O,
       N149_O,N150_O,N151_O,N152_O,N153_O,N154_O,N155_O,N156_O,N157_O,N158_O,
       N159_O,N160_O,N161_O,N162_O,N163_O,N164_O,N165_O,N166_O,N167_O,N168_O,
       N169_O,N170_O,N171_O,N172_O,N173_O,N174_O,N175_O,N176_O,N177_O,N178_O,
       N179_O,N180_O,N181_O,N182_O,N183_O,N184_O,N185_O,N186_O,N187_O,N188_O,
       N189_O,N190_O,N191_O,N192_O,N193_O,N194_O,N195_O,N196_O,N197_O,N198_O,
       N199_O,N200_O,N201_O,N202_O,N203_O,N204_O,N205_O,N206_O,N207_O,N208_O,
       N209_O,N210_O,N211_O,N212_O,N213_O,N214_O,N215_O,N216_O,N217_O,N218_O;

wire N405,N408,N425,N485,N486,N495,N496,N499,N500,N503,
     N506,N509,N521,N533,N537,N543,N544,N547,N550,N562,
     N574,N578,N582,N594,N606,N607,N608,N609,N610,N611,
     N612,N613,N625,N637,N643,N650,N651,N655,N659,N663,
     N667,N671,N675,N679,N683,N687,N693,N699,N705,N711,
     N715,N719,N723,N727,N730,N733,N734,N735,N738,N741,
     N744,N747,N750,N753,N756,N759,N762,N765,N768,N771,
     N774,N777,N780,N783,N786,N800,N900,N901,N902,N903,
     N904,N905,N998,N999,N1027,N1032,N1033,N1034,N1037,N1042,
     N1053,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1075,N1086,
     N1097,N1098,N1099,N1100,N1101,N1102,N1113,N1124,N1125,N1126,
     N1127,N1128,N1129,N1133,N1137,N1140,N1141,N1142,N1143,N1144,
     N1145,N1146,N1157,N1168,N1169,N1170,N1171,N1172,N1173,N1178,
     N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1195,N1200,N1205,
     N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1219,N1222,N1225,
     N1228,N1231,N1234,N1237,N1240,N1243,N1246,N1249,N1250,N1251,
     N1254,N1257,N1260,N1263,N1266,N1275,N1276,N1302,N1351,N1352,
     N1353,N1354,N1355,N1395,N1396,N1397,N1398,N1399,N1422,N1423,
     N1424,N1425,N1426,N1427,N1440,N1441,N1449,N1450,N1451,N1452,
     N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,
     N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,
     N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,
     N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,N1491,N1492,
     N1493,N1494,N1495,N1496,N1499,N1502,N1506,N1510,N1513,N1516,
     N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,
     N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,
     N1549,N1550,N1551,N1552,N1553,N1557,N1561,N1564,N1565,N1566,
     N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,
     N1577,N1578,N1581,N1582,N1585,N1588,N1591,N1596,N1600,N1606,
     N1612,N1615,N1619,N1624,N1628,N1631,N1634,N1637,N1642,N1647,
     N1651,N1656,N1676,N1681,N1686,N1690,N1708,N1770,N1773,N1776,
     N1777,N1778,N1781,N1784,N1785,N1795,N1798,N1801,N1804,N1807,
     N1808,N1809,N1810,N1811,N1813,N1814,N1815,N1822,N1823,N1824,
     N1827,N1830,N1831,N1832,N1833,N1836,N1841,N1848,N1852,N1856,
     N1863,N1870,N1875,N1880,N1885,N1888,N1891,N1894,N1897,N1908,
     N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,N1918,
     N1919,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,
     N1939,N1940,N1941,N1942,N1945,N1948,N1951,N1954,N1957,N1960,
     N1963,N1966,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2040,
     N2041,N2042,N2043,N2046,N2049,N2052,N2055,N2058,N2061,N2064,
     N2067,N2070,N2073,N2076,N2079,N2095,N2098,N2101,N2104,N2107,
     N2110,N2113,N2119,N2120,N2125,N2126,N2127,N2128,N2135,N2141,
     N2144,N2147,N2150,N2153,N2154,N2155,N2156,N2157,N2158,N2171,
     N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2185,N2188,N2191,
     N2194,N2197,N2200,N2201,N2204,N2207,N2210,N2213,N2216,N2219,
     N2234,N2235,N2236,N2237,N2250,N2266,N2269,N2291,N2294,N2297,
     N2298,N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,
     N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,N2318,
     N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,
     N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,
     N2339,N2340,N2354,N2355,N2356,N2357,N2358,N2359,N2364,N2365,
     N2366,N2367,N2368,N2372,N2373,N2374,N2375,N2376,N2377,N2382,
     N2386,N2391,N2395,N2400,N2403,N2406,N2407,N2408,N2409,N2410,
     N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2421,N2425,N2428,
     N2429,N2430,N2431,N2432,N2433,N2434,N2437,N2440,N2443,N2446,
     N2449,N2452,N2453,N2454,N2457,N2460,N2463,N2466,N2469,N2472,
     N2475,N2478,N2481,N2484,N2487,N2490,N2493,N2503,N2504,N2510,
     N2511,N2521,N2528,N2531,N2534,N2537,N2540,N2544,N2545,N2546,
     N2547,N2548,N2549,N2550,N2551,N2552,N2553,N2563,N2564,N2565,
     N2566,N2567,N2568,N2579,N2603,N2607,N2608,N2609,N2610,N2611,
     N2612,N2613,N2617,N2618,N2619,N2620,N2621,N2624,N2628,N2629,
     N2630,N2631,N2632,N2633,N2634,N2635,N2636,N2638,N2645,N2646,
     N2652,N2655,N2656,N2659,N2663,N2664,N2665,N2666,N2667,N2668,
     N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2677,N2678,
     N2679,N2680,N2681,N2684,N2687,N2690,N2693,N2694,N2695,N2696,
     N2697,N2698,N2699,N2700,N2701,N2702,N2703,N2706,N2707,N2708,
     N2709,N2710,N2719,N2720,N2726,N2729,N2738,N2743,N2747,N2748,
     N2749,N2750,N2751,N2760,N2761,N2766,N2771,N2772,N2773,N2774,
     N2775,N2776,N2777,N2778,N2781,N2782,N2783,N2784,N2789,N2790,
     N2791,N2792,N2793,N2796,N2800,N2803,N2806,N2809,N2810,N2811,
     N2812,N2817,N2820,N2826,N2829,N2830,N2831,N2837,N2838,N2839,
     N2840,N2841,N2844,N2854,N2859,N2869,N2874,N2877,N2880,N2881,
     N2882,N2885,N2888,N2894,N2895,N2896,N2897,N2898,N2899,N2900,
     N2901,N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2931,
     N2938,N2939,N2963,N2972,N2975,N2978,N2981,N2984,N2985,N2986,
     N2989,N2992,N2995,N2998,N3001,N3004,N3007,N3008,N3009,N3010,
     N3013,N3016,N3019,N3022,N3025,N3028,N3029,N3030,N3035,N3036,
     N3037,N3039,N3044,N3045,N3046,N3047,N3048,N3049,N3050,N3053,
     N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,N3064,N3065,
     N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,N3074,N3075,
     N3076,N3088,N3091,N3110,N3113,N3137,N3140,N3143,N3146,N3149,
     N3152,N3157,N3160,N3163,N3166,N3169,N3172,N3175,N3176,N3177,
     N3178,N3180,N3187,N3188,N3189,N3190,N3191,N3192,N3193,N3194,
     N3195,N3196,N3197,N3208,N3215,N3216,N3217,N3218,N3219,N3220,
     N3222,N3223,N3230,N3231,N3238,N3241,N3244,N3247,N3250,N3253,
     N3256,N3259,N3262,N3265,N3268,N3271,N3274,N3277,N3281,N3282,
     N3283,N3284,N3286,N3288,N3289,N3291,N3293,N3295,N3296,N3299,
     N3301,N3302,N3304,N3306,N3308,N3309,N3312,N3314,N3315,N3318,
     N3321,N3324,N3327,N3330,N3333,N3334,N3335,N3336,N3337,N3340,
     N3344,N3348,N3352,N3356,N3360,N3364,N3367,N3370,N3374,N3378,
     N3382,N3386,N3390,N3394,N3397,N3400,N3401,N3402,N3403,N3404,
     N3405,N3406,N3409,N3410,N3412,N3414,N3416,N3418,N3420,N3422,
     N3428,N3430,N3432,N3434,N3436,N3438,N3440,N3450,N3453,N3456,
     N3459,N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,N3486,
     N3487,N3488,N3489,N3490,N3491,N3492,N3493,N3494,N3496,N3498,
     N3499,N3500,N3501,N3502,N3503,N3504,N3505,N3506,N3507,N3508,
     N3509,N3510,N3511,N3512,N3513,N3515,N3517,N3522,N3525,N3528,
     N3531,N3534,N3537,N3540,N3543,N3551,N3552,N3553,N3554,N3555,
     N3556,N3557,N3558,N3559,N3563,N3564,N3565,N3566,N3567,N3568,
     N3569,N3570,N3576,N3579,N3585,N3588,N3592,N3593,N3594,N3595,
     N3596,N3597,N3598,N3599,N3600,N3603,N3608,N3612,N3615,N3616,
     N3622,N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3640,N3644,
     N3647,N3648,N3654,N3661,N3662,N3667,N3668,N3669,N3670,N3691,
     N3692,N3693,N3694,N3695,N3696,N3697,N3716,N3717,N3718,N3719,
     N3720,N3721,N3722,N3723,N3726,N3727,N3728,N3729,N3730,N3731,
     N3732,N3733,N3734,N3735,N3736,N3737,N3740,N3741,N3742,N3743,
     N3744,N3745,N3746,N3747,N3748,N3749,N3750,N3753,N3754,N3758,
     N3761,N3762,N3767,N3771,N3774,N3775,N3778,N3779,N3780,N3790,
     N3793,N3794,N3802,N3805,N3806,N3807,N3808,N3811,N3812,N3813,
     N3814,N3815,N3816,N3817,N3818,N3819,N3820,N3821,N3822,N3823,
     N3826,N3827,N3834,N3835,N3836,N3837,N3838,N3839,N3840,N3843,
     N3852,N3857,N3858,N3859,N3864,N3869,N3870,N3876,N3877,
     N11_NOT,N246_NOT,N7_NOT,N237_NOT,N343_NOT,N610_NOT,N340_NOT,N611_NOT,N547_NOT,N544_NOT,
     N904_NOT,N905_NOT,N744_NOT,N1143_NOT,N759_NOT,N1212_NOT,N1102_NOT,N594_NOT,N4_NOT,N1173_NOT,
     N22_NOT,N1178_NOT,N6_NOT,N1178_NOT,N1424_NOT,N1425_NOT,N1606_NOT,N241_NOT,N1606_NOT,N637_NOT,
     N1612_NOT,N637_NOT,N1619_NOT,N643_NOT,N1631_NOT,N643_NOT,N1634_NOT,N643_NOT,N1676_NOT,N693_NOT,
     N1637_NOT,N699_NOT,N1647_NOT,N699_NOT,N533_NOT,N1815_NOT,N1909_NOT,N1785_NOT,N1547_NOT,N1913_NOT,
     N1568_NOT,N1932_NOT,N1824_NOT,N537_NOT,N2157_NOT,N2032_NOT,N2052_NOT,N1519_NOT,N2055_NOT,N1520_NOT,
     N2076_NOT,N1527_NOT,N2098_NOT,N1573_NOT,N2110_NOT,N1577_NOT,N2120_NOT,N533_NOT,N1228_NOT,N2309_NOT,
     N1240_NOT,N2317_NOT,N1266_NOT,N2340_NOT,N2302_NOT,N2407_NOT,N2308_NOT,N2410_NOT,N2310_NOT,N2411_NOT,
     N2318_NOT,N2415_NOT,N1936_NOT,N2452_NOT,N1676_NOT,N2377_NOT,N1681_NOT,N2377_NOT,N1863_NOT,N2391_NOT,
     N1880_NOT,N2395_NOT,N2294_NOT,N2534_NOT,N2443_NOT,N2695_NOT,N2709_NOT,N2534_NOT,N1856_NOT,N2638_NOT,
     N2750_NOT,N2751_NOT,N2811_NOT,N1070_NOT,N2636_NOT,N2738_NOT,N578_NOT,N2831_NOT,N2938_NOT,N2839_NOT,
     N687_NOT,N2854_NOT,N663_NOT,N2859_NOT,N667_NOT,N2859_NOT,N679_NOT,N2869_NOT,N3056_NOT,N1190_NOT,
     N3059_NOT,N2761_NOT,N3066_NOT,N1195_NOT,N705_NOT,N3030_NOT,N719_NOT,N3050_NOT,N723_NOT,N3050_NOT,
     N719_NOT,N3061_NOT,N723_NOT,N3061_NOT,N2210_NOT,N3196_NOT,N3152_NOT,N2981_NOT,N3149_NOT,N2978_NOT,
     N3172_NOT,N3025_NOT,N3219_NOT,N3045_NOT,N3195_NOT,N3286_NOT,N3283_NOT,N3193_NOT,N3335_NOT,N1190_NOT,
     N3400_NOT,N533_NOT,N3315_NOT,N1841_NOT,N3344_NOT,N3414_NOT,N3370_NOT,N3430_NOT,N3378_NOT,N3434_NOT,
     N3404_NOT,N3403_NOT,N3250_NOT,N3486_NOT,N3528_NOT,N2630_NOT,N3531_NOT,N2376_NOT,N3554_NOT,N3487_NOT,
     N3555_NOT,N3489_NOT,N3556_NOT,N3491_NOT,N3537_NOT,N2655_NOT,N3564_NOT,N3504_NOT,N3238_NOT,N3592_NOT,
     N3576_NOT,N3494_NOT,N3729_NOT,N3694_NOT,N3737_NOT,N3500_NOT,N3816_NOT,N3817_NOT,N3818_NOT,N3823_NOT,
     EX1,EX2,EX3,EX4,EX5,EX6,EX7,EX8,EX9,EX10,
     EX11,EX12,EX13,EX14,EX15,EX16,EX17,EX18,EX19,EX20,
     EX21,EX22,EX23,EX24,EX25,EX26,EX27,EX28,EX29,EX30,
     EX31,EX32,EX33,EX34,EX35,EX36,EX37,EX38,EX39,EX40,
     EX41,EX42,EX43,EX44,EX45,EX46,EX47,EX48,EX49,EX50,
     EX51,EX52,EX53,EX54,EX55,EX56,EX57,EX58,EX59,EX60,
     EX61,EX62,EX63,EX64,EX65,EX66,EX67,EX68,EX69,EX70,
     EX71,EX72,EX73,EX74,EX75,EX76,EX77,EX78,EX79,EX80,
     EX81,EX82,EX83,EX84,EX85,EX86,EX87,EX88,EX89,EX90,
     EX91,EX92,EX93,EX94,EX95,EX96,EX97,EX98,EX99,EX100,
     EX101,EX102,EX103,EX104,EX105,EX106,EX107,EX108,EX109,EX110,
     EX111,EX112,EX113,EX114,EX115,EX116,EX117,EX118,EX119,EX120,
     EX121,EX122,EX123,EX124,EX125,EX126,EX127,EX128,EX129,EX130,
     EX131,EX132,EX133,EX134,EX135,EX136,EX137,EX138,EX139,EX140,
     EX141,EX142,EX143,EX144,EX145,EX146,EX147,EX148,EX149,EX150,
     EX151,EX152,EX153,EX154,EX155,EX156,EX157,EX158,EX159,EX160,
     EX161,EX162,EX163,EX164,EX165,EX166,EX167,EX168,EX169,EX170,
     EX171,EX172,EX173,EX174,EX175,EX176,EX177,EX178,EX179,EX180,
     EX181,EX182,EX183,EX184,EX185,EX186,EX187,EX188,EX189,EX190,
     EX191,EX192,EX193,EX194,EX195,EX196,EX197,EX198,EX199,EX200,
     EX201,EX202,EX203,EX204,EX205,EX206,EX207,EX208,EX209,EX210,
     EX211,EX212,EX213,EX214,EX215,EX216,EX217,EX218,EX219,EX220,
     EX221,EX222,EX223,EX224,EX225,EX226,EX227,EX228,EX229,EX230,
     EX231,EX232,EX233,EX234,EX235,EX236,EX237,EX238,EX239,EX240,
     EX241,EX242,EX243,EX244,EX245,EX246,EX247,EX248,EX249,EX250,
     EX251,EX252,EX253,EX254,EX255,EX256,EX257,EX258,EX259,EX260,
     EX261,EX262,EX263,EX264,EX265,EX266,EX267,EX268,EX269,EX270,
     EX271,EX272,EX273,EX274,EX275,EX276,EX277,EX278,EX279,EX280,
     EX281,EX282,EX283,EX284,EX285,EX286,EX287,EX288,EX289,EX290,
     EX291,EX292,EX293,EX294,EX295,EX296,EX297,EX298,EX299,EX300,
     EX301,EX302,EX303,EX304,EX305,EX306,EX307,EX308,EX309,EX310,
     EX311,EX312,EX313,EX314,EX315,EX316,EX317,EX318,EX319,EX320,
     EX321,EX322,EX323,EX324,EX325,EX326,EX327,EX328,EX329,EX330,
     EX331,EX332,EX333,EX334,EX335,EX336,EX337,EX338,EX339,EX340,
     EX341,EX342,EX343,EX344,EX345,EX346,EX347,EX348,EX349,EX350,
     EX351,EX352,EX353,EX354,EX355,EX356,EX357,EX358,EX359,EX360,
     EX361,EX362,EX363,EX364,EX365,EX366,EX367,EX368,EX369,EX370,
     EX371,EX372,EX373,EX374,EX375,EX376,EX377,EX378,EX379,EX380,
     EX381,EX382,EX383,EX384,EX385,EX386,EX387,EX388,EX389,EX390,
     EX391,EX392,EX393,EX394,EX395,EX396,EX397,EX398,EX399,EX400,
     EX401,EX402,EX403,EX404,EX405,EX406,EX407,EX408,EX409,EX410,
     EX411,EX412,EX413,EX414,EX415,EX416,EX417,EX418,EX419,EX420,
     EX421,EX422,EX423,EX424,EX425,EX426,EX427,EX428,EX429,EX430,
     EX431,EX432,EX433,EX434,EX435,EX436,EX437,EX438,EX439,EX440,
     EX441,EX442,EX443,EX444,EX445,EX446,EX447,EX448,EX449,EX450,
     EX451,EX452,EX453,EX454,EX455,EX456,EX457,EX458,EX459,EX460,
     EX461,EX462,EX463,EX464,EX465,EX466,EX467,EX468,EX469,EX470,
     EX471,EX472,EX473,EX474,EX475,EX476,EX477,EX478,EX479,EX480,
     EX481,EX482,EX483,EX484,EX485,EX486,EX487,EX488,EX489,EX490,
     EX491,EX492,EX493,EX494,EX495,EX496,EX497,EX498,EX499,EX500,
     EX501,EX502,EX503,EX504,EX505,EX506,EX507,EX508,EX509,EX510,
     EX511,EX512,EX513,EX514,EX515,EX516,EX517,EX518,EX519,EX520,
     EX521,EX522,EX523,EX524,EX525,EX526,EX527,EX528,EX529,EX530,
     EX531,EX532,EX533,EX534,EX535,EX536,EX537,EX538,EX539,EX540,
     EX541,EX542,EX543,EX544,EX545,EX546,EX547,EX548,EX549,EX550,
     EX551,EX552,EX553,EX554,EX555,EX556,EX557,EX558,EX559,EX560,
     EX561,EX562,EX563,EX564,EX565,EX566,EX567,EX568,EX569,EX570,
     EX571,EX572,EX573,EX574,EX575,EX576,EX577,EX578,EX579,EX580,
     EX581,EX582,EX583,EX584,EX585,EX586,EX587,EX588,EX589,EX590,
     EX591,EX592,EX593,EX594,EX595,EX596,EX597,EX598,EX599,EX600,
     EX601,EX602,EX603,EX604,EX605,EX606,EX607,EX608,EX609,EX610,
     EX611,EX612,EX613,EX614,EX615,EX616,EX617,EX618,EX619,EX620,
     EX621,EX622,EX623,EX624,EX625,EX626,EX627,EX628,EX629,EX630,
     EX631,EX632,EX633,EX634,EX635,EX636,EX637,EX638,EX639,EX640,
     EX641,EX642,EX643,EX644,EX645,EX646,EX647,EX648,EX649,EX650,
     EX651,EX652,EX653,EX654,EX655,EX656,EX657,EX658,EX659,EX660,
     EX661,EX662,EX663,EX664,EX665,EX666,EX667,EX668,EX669,EX670,
     EX671,EX672,EX673,EX674,EX675,EX676,EX677,EX678,EX679,EX680,
     EX681,EX682,EX683,EX684,EX685,EX686,EX687,EX688,EX689,EX690,
     EX691,EX692,EX693,EX694,EX695,EX696,EX697,EX698,EX699,EX700,
     EX701,EX702,EX703,EX704,EX705,EX706,EX707,EX708,EX709,EX710,
     EX711,EX712,EX713,EX714,EX715,EX716,EX717,EX718,EX719,EX720,
     EX721,EX722,EX723,EX724,EX725,EX726,EX727,EX728,EX729,EX730,
     EX731,EX732,EX733,EX734,EX735,EX736,EX737,EX738,EX739,EX740,
     EX741,EX742,EX743,EX744,EX745,EX746,EX747,EX748,EX749,EX750,
     EX751,EX752,EX753,EX754,EX755,EX756,EX757,EX758,EX759,EX760,
     EX761,EX762,EX763,EX764,EX765,EX766,EX767,EX768,EX769,EX770,
     EX771,EX772,EX773,EX774,EX775,EX776,EX777,EX778,EX779,EX780,
     EX781,EX782,EX783,EX784,EX785,EX786,EX787,EX788,EX789,EX790,
     EX791,EX792,EX793,EX794,EX795,EX796,EX797,EX798,EX799,EX800,
     EX801,EX802,EX803,EX804,EX805,EX806,EX807,EX808,EX809,EX810,
     EX811,EX812,EX813,EX814,EX815,EX816,EX817,EX818,EX819,EX820,
     EX821,EX822,EX823,EX824,EX825,EX826,EX827,EX828,EX829,EX830,
     EX831,EX832,EX833,EX834,EX835,EX836,EX837,EX838,EX839,EX840,
     EX841,EX842,EX843,EX844,EX845,EX846,EX847,EX848,EX849,EX850,
     EX851,EX852,EX853,EX854,EX855,EX856,EX857,EX858,EX859,EX860,
     EX861,EX862,EX863,EX864,EX865,EX866,EX867,EX868,EX869,EX870,
     EX871,EX872,EX873,EX874,EX875,EX876,EX877,EX878,EX879,EX880,
     EX881,EX882,EX883,EX884,EX885,EX886,EX887,EX888,EX889,EX890,
     EX891,EX892,EX893,EX894,EX895,EX896,EX897,EX898,EX899,EX900,
     EX901,EX902,EX903,EX904,EX905,EX906,EX907,EX908,EX909,EX910,
     EX911,EX912,EX913,EX914,EX915,EX916,EX917,EX918,EX919,EX920,
     EX921,EX922,EX923,EX924,EX925,EX926,EX927,EX928,EX929,EX930,
     EX931,EX932,EX933,EX934,EX935,EX936,EX937,EX938,EX939,EX940,
     EX941,EX942,EX943,EX944,EX945,EX946,EX947,EX948,EX949,EX950;


buf1 gate1( .a(N219), .O(N398) );
buf1 gate2( .a(N219), .O(N400) );
buf1 gate3( .a(N219), .O(N401) );
and2 gate4( .a(N1), .b(N3), .O(N405) );
inv1 gate5( .a(N230), .O(N408) );
buf1 gate6( .a(N253), .O(N419) );
buf1 gate7( .a(N253), .O(N420) );
inv1 gate8( .a(N262), .O(N425) );
buf1 gate9( .a(N290), .O(N456) );
buf1 gate10( .a(N290), .O(N457) );
buf1 gate11( .a(N290), .O(N458) );
and4 gate12( .a(N309), .b(N305), .c(N301), .d(N297), .O(N485) );
inv1 gate13( .a(N405), .O(N486) );
inv1 gate14( .a(N44), .O(N487) );
inv1 gate15( .a(N132), .O(N488) );
inv1 gate16( .a(N82), .O(N489) );
inv1 gate17( .a(N96), .O(N490) );
inv1 gate18( .a(N69), .O(N491) );
inv1 gate19( .a(N120), .O(N492) );
inv1 gate20( .a(N57), .O(N493) );
inv1 gate21( .a(N108), .O(N494) );
and3 gate22( .a(N2), .b(N15), .c(N237), .O(N495) );
buf1 gate23( .a(N237), .O(N496) );
and2 gate24( .a(N37), .b(N37), .O(N499) );
buf1 gate25( .a(N219), .O(N500) );
buf1 gate26( .a(N8), .O(N503) );
buf1 gate27( .a(N8), .O(N506) );
buf1 gate28( .a(N227), .O(N509) );
buf1 gate29( .a(N234), .O(N521) );
inv1 gate30( .a(N241), .O(N533) );
inv1 gate31( .a(N246), .O(N537) );
inv1 gate( .a(N11),.O(N11_NOT) );
inv1 gate( .a(N246),.O(N246_NOT));
and2 gate( .a(N11_NOT), .b(p1), .O(EX1) );
and2 gate( .a(N246_NOT), .b(EX1), .O(EX2) );
and2 gate( .a(N11), .b(p2), .O(EX3) );
and2 gate( .a(N246_NOT), .b(EX3), .O(EX4) );
and2 gate( .a(N11_NOT), .b(p3), .O(EX5) );
and2 gate( .a(N246), .b(EX5), .O(EX6) );
and2 gate( .a(N11), .b(p4), .O(EX7) );
and2 gate( .a(N246), .b(EX7), .O(EX8) );
or2  gate( .a(EX2), .b(EX4), .O(EX9) );
or2  gate( .a(EX6), .b(EX9), .O(EX10) );
or2  gate( .a(EX8), .b(EX10), .O(N543) );
and4 gate33( .a(N132), .b(N82), .c(N96), .d(N44), .O(N544) );
and4 gate34( .a(N120), .b(N57), .c(N108), .d(N69), .O(N547) );
buf1 gate35( .a(N227), .O(N550) );
buf1 gate36( .a(N234), .O(N562) );
inv1 gate37( .a(N256), .O(N574) );
inv1 gate38( .a(N259), .O(N578) );
buf1 gate39( .a(N319), .O(N582) );
buf1 gate40( .a(N322), .O(N594) );
inv1 gate41( .a(N328), .O(N606) );
inv1 gate42( .a(N331), .O(N607) );
inv1 gate43( .a(N334), .O(N608) );
inv1 gate44( .a(N337), .O(N609) );
inv1 gate45( .a(N340), .O(N610) );
inv1 gate46( .a(N343), .O(N611) );
inv1 gate47( .a(N352), .O(N612) );
buf1 gate48( .a(N319), .O(N613) );
buf1 gate49( .a(N322), .O(N625) );
buf1 gate50( .a(N16), .O(N637) );
buf1 gate51( .a(N16), .O(N643) );
inv1 gate52( .a(N355), .O(N650) );
inv1 gate( .a(N7),.O(N7_NOT) );
inv1 gate( .a(N237),.O(N237_NOT));
and2 gate( .a(N7_NOT), .b(p5), .O(EX11) );
and2 gate( .a(N237_NOT), .b(EX11), .O(EX12) );
and2 gate( .a(N7), .b(p6), .O(EX13) );
and2 gate( .a(N237_NOT), .b(EX13), .O(EX14) );
and2 gate( .a(N7_NOT), .b(p7), .O(EX15) );
and2 gate( .a(N237), .b(EX15), .O(EX16) );
and2 gate( .a(N7), .b(p8), .O(EX17) );
and2 gate( .a(N237), .b(EX17), .O(EX18) );
or2  gate( .a(EX12), .b(EX14), .O(EX19) );
or2  gate( .a(EX16), .b(EX19), .O(EX20) );
or2  gate( .a(EX18), .b(EX20), .O(N651) );
inv1 gate54( .a(N263), .O(N655) );
inv1 gate55( .a(N266), .O(N659) );
inv1 gate56( .a(N269), .O(N663) );
inv1 gate57( .a(N272), .O(N667) );
inv1 gate58( .a(N275), .O(N671) );
inv1 gate59( .a(N278), .O(N675) );
inv1 gate60( .a(N281), .O(N679) );
inv1 gate61( .a(N284), .O(N683) );
inv1 gate62( .a(N287), .O(N687) );
buf1 gate63( .a(N29), .O(N693) );
buf1 gate64( .a(N29), .O(N699) );
inv1 gate65( .a(N294), .O(N705) );
inv1 gate66( .a(N297), .O(N711) );
inv1 gate67( .a(N301), .O(N715) );
inv1 gate68( .a(N305), .O(N719) );
inv1 gate69( .a(N309), .O(N723) );
inv1 gate70( .a(N313), .O(N727) );
inv1 gate71( .a(N316), .O(N730) );
inv1 gate72( .a(N346), .O(N733) );
inv1 gate73( .a(N349), .O(N734) );
buf1 gate74( .a(N259), .O(N735) );
buf1 gate75( .a(N256), .O(N738) );
buf1 gate76( .a(N263), .O(N741) );
buf1 gate77( .a(N269), .O(N744) );
buf1 gate78( .a(N266), .O(N747) );
buf1 gate79( .a(N275), .O(N750) );
buf1 gate80( .a(N272), .O(N753) );
buf1 gate81( .a(N281), .O(N756) );
buf1 gate82( .a(N278), .O(N759) );
buf1 gate83( .a(N287), .O(N762) );
buf1 gate84( .a(N284), .O(N765) );
buf1 gate85( .a(N294), .O(N768) );
buf1 gate86( .a(N301), .O(N771) );
buf1 gate87( .a(N297), .O(N774) );
buf1 gate88( .a(N309), .O(N777) );
buf1 gate89( .a(N305), .O(N780) );
buf1 gate90( .a(N316), .O(N783) );
buf1 gate91( .a(N313), .O(N786) );
inv1 gate92( .a(N485), .O(N792) );
inv1 gate93( .a(N495), .O(N799) );
inv1 gate94( .a(N499), .O(N800) );
buf1 gate95( .a(N500), .O(N805) );
nand2 gate96( .a(N331), .b(N606), .O(N900) );
nand2 gate97( .a(N328), .b(N607), .O(N901) );
nand2 gate98( .a(N337), .b(N608), .O(N902) );
nand2 gate99( .a(N334), .b(N609), .O(N903) );
inv1 gate( .a(N343),.O(N343_NOT) );
inv1 gate( .a(N610),.O(N610_NOT));
and2 gate( .a(N343_NOT), .b(p9), .O(EX21) );
and2 gate( .a(N610_NOT), .b(EX21), .O(EX22) );
and2 gate( .a(N343), .b(p10), .O(EX23) );
and2 gate( .a(N610_NOT), .b(EX23), .O(EX24) );
and2 gate( .a(N343_NOT), .b(p11), .O(EX25) );
and2 gate( .a(N610), .b(EX25), .O(EX26) );
and2 gate( .a(N343), .b(p12), .O(EX27) );
and2 gate( .a(N610), .b(EX27), .O(EX28) );
or2  gate( .a(EX22), .b(EX24), .O(EX29) );
or2  gate( .a(EX26), .b(EX29), .O(EX30) );
or2  gate( .a(EX28), .b(EX30), .O(N904) );
inv1 gate( .a(N340),.O(N340_NOT) );
inv1 gate( .a(N611),.O(N611_NOT));
and2 gate( .a(N340_NOT), .b(p13), .O(EX31) );
and2 gate( .a(N611_NOT), .b(EX31), .O(EX32) );
and2 gate( .a(N340), .b(p14), .O(EX33) );
and2 gate( .a(N611_NOT), .b(EX33), .O(EX34) );
and2 gate( .a(N340_NOT), .b(p15), .O(EX35) );
and2 gate( .a(N611), .b(EX35), .O(EX36) );
and2 gate( .a(N340), .b(p16), .O(EX37) );
and2 gate( .a(N611), .b(EX37), .O(EX38) );
or2  gate( .a(EX32), .b(EX34), .O(EX39) );
or2  gate( .a(EX36), .b(EX39), .O(EX40) );
or2  gate( .a(EX38), .b(EX40), .O(N905) );
nand2 gate102( .a(N349), .b(N733), .O(N998) );
nand2 gate103( .a(N346), .b(N734), .O(N999) );
and2 gate104( .a(N94), .b(N500), .O(N1026) );
and2 gate105( .a(N325), .b(N651), .O(N1027) );
inv1 gate106( .a(N651), .O(N1028) );
nand2 gate107( .a(N231), .b(N651), .O(N1029) );
inv1 gate108( .a(N544), .O(N1032) );
inv1 gate109( .a(N547), .O(N1033) );
inv1 gate( .a(N547),.O(N547_NOT) );
inv1 gate( .a(N544),.O(N544_NOT));
and2 gate( .a(N547_NOT), .b(p17), .O(EX41) );
and2 gate( .a(N544_NOT), .b(EX41), .O(EX42) );
and2 gate( .a(N547), .b(p18), .O(EX43) );
and2 gate( .a(N544_NOT), .b(EX43), .O(EX44) );
and2 gate( .a(N547_NOT), .b(p19), .O(EX45) );
and2 gate( .a(N544), .b(EX45), .O(EX46) );
and2 gate( .a(N547), .b(p20), .O(EX47) );
and2 gate( .a(N544), .b(EX47), .O(EX48) );
or2  gate( .a(EX42), .b(EX44), .O(EX49) );
or2  gate( .a(EX46), .b(EX49), .O(EX50) );
or2  gate( .a(EX48), .b(EX50), .O(N1034) );
buf1 gate111( .a(N503), .O(N1037) );
inv1 gate112( .a(N509), .O(N1042) );
inv1 gate113( .a(N521), .O(N1053) );
and3 gate114( .a(N80), .b(N509), .c(N521), .O(N1064) );
and3 gate115( .a(N68), .b(N509), .c(N521), .O(N1065) );
and3 gate116( .a(N79), .b(N509), .c(N521), .O(N1066) );
and3 gate117( .a(N78), .b(N509), .c(N521), .O(N1067) );
and3 gate118( .a(N77), .b(N509), .c(N521), .O(N1068) );
and2 gate119( .a(N11), .b(N537), .O(N1069) );
buf1 gate120( .a(N503), .O(N1070) );
inv1 gate121( .a(N550), .O(N1075) );
inv1 gate122( .a(N562), .O(N1086) );
and3 gate123( .a(N76), .b(N550), .c(N562), .O(N1097) );
and3 gate124( .a(N75), .b(N550), .c(N562), .O(N1098) );
and3 gate125( .a(N74), .b(N550), .c(N562), .O(N1099) );
and3 gate126( .a(N73), .b(N550), .c(N562), .O(N1100) );
and3 gate127( .a(N72), .b(N550), .c(N562), .O(N1101) );
inv1 gate128( .a(N582), .O(N1102) );
inv1 gate129( .a(N594), .O(N1113) );
and3 gate130( .a(N114), .b(N582), .c(N594), .O(N1124) );
and3 gate131( .a(N113), .b(N582), .c(N594), .O(N1125) );
and3 gate132( .a(N112), .b(N582), .c(N594), .O(N1126) );
and3 gate133( .a(N111), .b(N582), .c(N594), .O(N1127) );
and2 gate134( .a(N582), .b(N594), .O(N1128) );
nand2 gate135( .a(N900), .b(N901), .O(N1129) );
nand2 gate136( .a(N902), .b(N903), .O(N1133) );
inv1 gate( .a(N904),.O(N904_NOT) );
inv1 gate( .a(N905),.O(N905_NOT));
and2 gate( .a(N904_NOT), .b(p21), .O(EX51) );
and2 gate( .a(N905_NOT), .b(EX51), .O(EX52) );
and2 gate( .a(N904), .b(p22), .O(EX53) );
and2 gate( .a(N905_NOT), .b(EX53), .O(EX54) );
and2 gate( .a(N904_NOT), .b(p23), .O(EX55) );
and2 gate( .a(N905), .b(EX55), .O(EX56) );
and2 gate( .a(N904), .b(p24), .O(EX57) );
and2 gate( .a(N905), .b(EX57), .O(EX58) );
or2  gate( .a(EX52), .b(EX54), .O(EX59) );
or2  gate( .a(EX56), .b(EX59), .O(EX60) );
or2  gate( .a(EX58), .b(EX60), .O(N1137) );
inv1 gate138( .a(N741), .O(N1140) );
nand2 gate139( .a(N741), .b(N612), .O(N1141) );
inv1 gate140( .a(N744), .O(N1142) );
inv1 gate141( .a(N747), .O(N1143) );
inv1 gate142( .a(N750), .O(N1144) );
inv1 gate143( .a(N753), .O(N1145) );
inv1 gate144( .a(N613), .O(N1146) );
inv1 gate145( .a(N625), .O(N1157) );
and3 gate146( .a(N118), .b(N613), .c(N625), .O(N1168) );
and3 gate147( .a(N107), .b(N613), .c(N625), .O(N1169) );
and3 gate148( .a(N117), .b(N613), .c(N625), .O(N1170) );
and3 gate149( .a(N116), .b(N613), .c(N625), .O(N1171) );
and3 gate150( .a(N115), .b(N613), .c(N625), .O(N1172) );
inv1 gate151( .a(N637), .O(N1173) );
inv1 gate152( .a(N643), .O(N1178) );
inv1 gate153( .a(N768), .O(N1184) );
nand2 gate154( .a(N768), .b(N650), .O(N1185) );
inv1 gate155( .a(N771), .O(N1186) );
inv1 gate156( .a(N774), .O(N1187) );
inv1 gate157( .a(N777), .O(N1188) );
inv1 gate158( .a(N780), .O(N1189) );
buf1 gate159( .a(N506), .O(N1190) );
buf1 gate160( .a(N506), .O(N1195) );
inv1 gate161( .a(N693), .O(N1200) );
inv1 gate162( .a(N699), .O(N1205) );
inv1 gate163( .a(N735), .O(N1210) );
inv1 gate164( .a(N738), .O(N1211) );
inv1 gate165( .a(N756), .O(N1212) );
inv1 gate166( .a(N759), .O(N1213) );
inv1 gate167( .a(N762), .O(N1214) );
inv1 gate168( .a(N765), .O(N1215) );
nand2 gate169( .a(N998), .b(N999), .O(N1216) );
buf1 gate170( .a(N574), .O(N1219) );
buf1 gate171( .a(N578), .O(N1222) );
buf1 gate172( .a(N655), .O(N1225) );
buf1 gate173( .a(N659), .O(N1228) );
buf1 gate174( .a(N663), .O(N1231) );
buf1 gate175( .a(N667), .O(N1234) );
buf1 gate176( .a(N671), .O(N1237) );
buf1 gate177( .a(N675), .O(N1240) );
buf1 gate178( .a(N679), .O(N1243) );
buf1 gate179( .a(N683), .O(N1246) );
inv1 gate180( .a(N783), .O(N1249) );
inv1 gate181( .a(N786), .O(N1250) );
buf1 gate182( .a(N687), .O(N1251) );
buf1 gate183( .a(N705), .O(N1254) );
buf1 gate184( .a(N711), .O(N1257) );
buf1 gate185( .a(N715), .O(N1260) );
buf1 gate186( .a(N719), .O(N1263) );
buf1 gate187( .a(N723), .O(N1266) );
inv1 gate188( .a(N1027), .O(N1269) );
and2 gate189( .a(N325), .b(N1032), .O(N1275) );
and2 gate190( .a(N231), .b(N1033), .O(N1276) );
buf1 gate191( .a(N1034), .O(N1277) );
or2 gate192( .a(N1069), .b(N543), .O(N1302) );
nand2 gate193( .a(N352), .b(N1140), .O(N1351) );
nand2 gate194( .a(N747), .b(N1142), .O(N1352) );
inv1 gate( .a(N744),.O(N744_NOT) );
inv1 gate( .a(N1143),.O(N1143_NOT));
and2 gate( .a(N744_NOT), .b(p25), .O(EX61) );
and2 gate( .a(N1143_NOT), .b(EX61), .O(EX62) );
and2 gate( .a(N744), .b(p26), .O(EX63) );
and2 gate( .a(N1143_NOT), .b(EX63), .O(EX64) );
and2 gate( .a(N744_NOT), .b(p27), .O(EX65) );
and2 gate( .a(N1143), .b(EX65), .O(EX66) );
and2 gate( .a(N744), .b(p28), .O(EX67) );
and2 gate( .a(N1143), .b(EX67), .O(EX68) );
or2  gate( .a(EX62), .b(EX64), .O(EX69) );
or2  gate( .a(EX66), .b(EX69), .O(EX70) );
or2  gate( .a(EX68), .b(EX70), .O(N1353) );
nand2 gate196( .a(N753), .b(N1144), .O(N1354) );
nand2 gate197( .a(N750), .b(N1145), .O(N1355) );
nand2 gate198( .a(N355), .b(N1184), .O(N1395) );
nand2 gate199( .a(N774), .b(N1186), .O(N1396) );
nand2 gate200( .a(N771), .b(N1187), .O(N1397) );
nand2 gate201( .a(N780), .b(N1188), .O(N1398) );
nand2 gate202( .a(N777), .b(N1189), .O(N1399) );
nand2 gate203( .a(N738), .b(N1210), .O(N1422) );
nand2 gate204( .a(N735), .b(N1211), .O(N1423) );
inv1 gate( .a(N759),.O(N759_NOT) );
inv1 gate( .a(N1212),.O(N1212_NOT));
and2 gate( .a(N759_NOT), .b(p29), .O(EX71) );
and2 gate( .a(N1212_NOT), .b(EX71), .O(EX72) );
and2 gate( .a(N759), .b(p30), .O(EX73) );
and2 gate( .a(N1212_NOT), .b(EX73), .O(EX74) );
and2 gate( .a(N759_NOT), .b(p31), .O(EX75) );
and2 gate( .a(N1212), .b(EX75), .O(EX76) );
and2 gate( .a(N759), .b(p32), .O(EX77) );
and2 gate( .a(N1212), .b(EX77), .O(EX78) );
or2  gate( .a(EX72), .b(EX74), .O(EX79) );
or2  gate( .a(EX76), .b(EX79), .O(EX80) );
or2  gate( .a(EX78), .b(EX80), .O(N1424) );
nand2 gate206( .a(N756), .b(N1213), .O(N1425) );
nand2 gate207( .a(N765), .b(N1214), .O(N1426) );
nand2 gate208( .a(N762), .b(N1215), .O(N1427) );
nand2 gate209( .a(N786), .b(N1249), .O(N1440) );
nand2 gate210( .a(N783), .b(N1250), .O(N1441) );
inv1 gate211( .a(N1034), .O(N1448) );
inv1 gate212( .a(N1275), .O(N1449) );
inv1 gate213( .a(N1276), .O(N1450) );
and3 gate214( .a(N93), .b(N1042), .c(N1053), .O(N1451) );
and3 gate215( .a(N55), .b(N509), .c(N1053), .O(N1452) );
and3 gate216( .a(N67), .b(N1042), .c(N521), .O(N1453) );
and3 gate217( .a(N81), .b(N1042), .c(N1053), .O(N1454) );
and3 gate218( .a(N43), .b(N509), .c(N1053), .O(N1455) );
and3 gate219( .a(N56), .b(N1042), .c(N521), .O(N1456) );
and3 gate220( .a(N92), .b(N1042), .c(N1053), .O(N1457) );
and3 gate221( .a(N54), .b(N509), .c(N1053), .O(N1458) );
and3 gate222( .a(N66), .b(N1042), .c(N521), .O(N1459) );
and3 gate223( .a(N91), .b(N1042), .c(N1053), .O(N1460) );
and3 gate224( .a(N53), .b(N509), .c(N1053), .O(N1461) );
and3 gate225( .a(N65), .b(N1042), .c(N521), .O(N1462) );
and3 gate226( .a(N90), .b(N1042), .c(N1053), .O(N1463) );
and3 gate227( .a(N52), .b(N509), .c(N1053), .O(N1464) );
and3 gate228( .a(N64), .b(N1042), .c(N521), .O(N1465) );
and3 gate229( .a(N89), .b(N1075), .c(N1086), .O(N1466) );
and3 gate230( .a(N51), .b(N550), .c(N1086), .O(N1467) );
and3 gate231( .a(N63), .b(N1075), .c(N562), .O(N1468) );
and3 gate232( .a(N88), .b(N1075), .c(N1086), .O(N1469) );
and3 gate233( .a(N50), .b(N550), .c(N1086), .O(N1470) );
and3 gate234( .a(N62), .b(N1075), .c(N562), .O(N1471) );
and3 gate235( .a(N87), .b(N1075), .c(N1086), .O(N1472) );
and3 gate236( .a(N49), .b(N550), .c(N1086), .O(N1473) );
and2 gate237( .a(N1075), .b(N562), .O(N1474) );
and3 gate238( .a(N86), .b(N1075), .c(N1086), .O(N1475) );
and3 gate239( .a(N48), .b(N550), .c(N1086), .O(N1476) );
and3 gate240( .a(N61), .b(N1075), .c(N562), .O(N1477) );
and3 gate241( .a(N85), .b(N1075), .c(N1086), .O(N1478) );
and3 gate242( .a(N47), .b(N550), .c(N1086), .O(N1479) );
and3 gate243( .a(N60), .b(N1075), .c(N562), .O(N1480) );
and3 gate244( .a(N138), .b(N1102), .c(N1113), .O(N1481) );
and3 gate245( .a(N102), .b(N582), .c(N1113), .O(N1482) );
and3 gate246( .a(N126), .b(N1102), .c(N594), .O(N1483) );
and3 gate247( .a(N137), .b(N1102), .c(N1113), .O(N1484) );
and3 gate248( .a(N101), .b(N582), .c(N1113), .O(N1485) );
and3 gate249( .a(N125), .b(N1102), .c(N594), .O(N1486) );
and3 gate250( .a(N136), .b(N1102), .c(N1113), .O(N1487) );
and3 gate251( .a(N100), .b(N582), .c(N1113), .O(N1488) );
and3 gate252( .a(N124), .b(N1102), .c(N594), .O(N1489) );
and3 gate253( .a(N135), .b(N1102), .c(N1113), .O(N1490) );
and3 gate254( .a(N99), .b(N582), .c(N1113), .O(N1491) );
and3 gate255( .a(N123), .b(N1102), .c(N594), .O(N1492) );
and2 gate256( .a(N1102), .b(N1113), .O(N1493) );
and2 gate257( .a(N582), .b(N1113), .O(N1494) );
inv1 gate( .a(N1102),.O(N1102_NOT) );
inv1 gate( .a(N594),.O(N594_NOT));
and2 gate( .a(N1102_NOT), .b(p33), .O(EX81) );
and2 gate( .a(N594_NOT), .b(EX81), .O(EX82) );
and2 gate( .a(N1102), .b(p34), .O(EX83) );
and2 gate( .a(N594_NOT), .b(EX83), .O(EX84) );
and2 gate( .a(N1102_NOT), .b(p35), .O(EX85) );
and2 gate( .a(N594), .b(EX85), .O(EX86) );
and2 gate( .a(N1102), .b(p36), .O(EX87) );
and2 gate( .a(N594), .b(EX87), .O(EX88) );
or2  gate( .a(EX82), .b(EX84), .O(EX89) );
or2  gate( .a(EX86), .b(EX89), .O(EX90) );
or2  gate( .a(EX88), .b(EX90), .O(N1495) );
inv1 gate259( .a(N1129), .O(N1496) );
inv1 gate260( .a(N1133), .O(N1499) );
nand2 gate261( .a(N1351), .b(N1141), .O(N1502) );
nand2 gate262( .a(N1352), .b(N1353), .O(N1506) );
nand2 gate263( .a(N1354), .b(N1355), .O(N1510) );
buf1 gate264( .a(N1137), .O(N1513) );
buf1 gate265( .a(N1137), .O(N1516) );
inv1 gate266( .a(N1219), .O(N1519) );
inv1 gate267( .a(N1222), .O(N1520) );
inv1 gate268( .a(N1225), .O(N1521) );
inv1 gate269( .a(N1228), .O(N1522) );
inv1 gate270( .a(N1231), .O(N1523) );
inv1 gate271( .a(N1234), .O(N1524) );
inv1 gate272( .a(N1237), .O(N1525) );
inv1 gate273( .a(N1240), .O(N1526) );
inv1 gate274( .a(N1243), .O(N1527) );
inv1 gate275( .a(N1246), .O(N1528) );
and3 gate276( .a(N142), .b(N1146), .c(N1157), .O(N1529) );
and3 gate277( .a(N106), .b(N613), .c(N1157), .O(N1530) );
and3 gate278( .a(N130), .b(N1146), .c(N625), .O(N1531) );
and3 gate279( .a(N131), .b(N1146), .c(N1157), .O(N1532) );
and3 gate280( .a(N95), .b(N613), .c(N1157), .O(N1533) );
and3 gate281( .a(N119), .b(N1146), .c(N625), .O(N1534) );
and3 gate282( .a(N141), .b(N1146), .c(N1157), .O(N1535) );
and3 gate283( .a(N105), .b(N613), .c(N1157), .O(N1536) );
and3 gate284( .a(N129), .b(N1146), .c(N625), .O(N1537) );
and3 gate285( .a(N140), .b(N1146), .c(N1157), .O(N1538) );
and3 gate286( .a(N104), .b(N613), .c(N1157), .O(N1539) );
and3 gate287( .a(N128), .b(N1146), .c(N625), .O(N1540) );
and3 gate288( .a(N139), .b(N1146), .c(N1157), .O(N1541) );
and3 gate289( .a(N103), .b(N613), .c(N1157), .O(N1542) );
and3 gate290( .a(N127), .b(N1146), .c(N625), .O(N1543) );
and2 gate291( .a(N19), .b(N1173), .O(N1544) );
inv1 gate( .a(N4),.O(N4_NOT) );
inv1 gate( .a(N1173),.O(N1173_NOT));
and2 gate( .a(N4_NOT), .b(p37), .O(EX91) );
and2 gate( .a(N1173_NOT), .b(EX91), .O(EX92) );
and2 gate( .a(N4), .b(p38), .O(EX93) );
and2 gate( .a(N1173_NOT), .b(EX93), .O(EX94) );
and2 gate( .a(N4_NOT), .b(p39), .O(EX95) );
and2 gate( .a(N1173), .b(EX95), .O(EX96) );
and2 gate( .a(N4), .b(p40), .O(EX97) );
and2 gate( .a(N1173), .b(EX97), .O(EX98) );
or2  gate( .a(EX92), .b(EX94), .O(EX99) );
or2  gate( .a(EX96), .b(EX99), .O(EX100) );
or2  gate( .a(EX98), .b(EX100), .O(N1545) );
and2 gate293( .a(N20), .b(N1173), .O(N1546) );
and2 gate294( .a(N5), .b(N1173), .O(N1547) );
and2 gate295( .a(N21), .b(N1178), .O(N1548) );
inv1 gate( .a(N22),.O(N22_NOT) );
inv1 gate( .a(N1178),.O(N1178_NOT));
and2 gate( .a(N22_NOT), .b(p41), .O(EX101) );
and2 gate( .a(N1178_NOT), .b(EX101), .O(EX102) );
and2 gate( .a(N22), .b(p42), .O(EX103) );
and2 gate( .a(N1178_NOT), .b(EX103), .O(EX104) );
and2 gate( .a(N22_NOT), .b(p43), .O(EX105) );
and2 gate( .a(N1178), .b(EX105), .O(EX106) );
and2 gate( .a(N22), .b(p44), .O(EX107) );
and2 gate( .a(N1178), .b(EX107), .O(EX108) );
or2  gate( .a(EX102), .b(EX104), .O(EX109) );
or2  gate( .a(EX106), .b(EX109), .O(EX110) );
or2  gate( .a(EX108), .b(EX110), .O(N1549) );
and2 gate297( .a(N23), .b(N1178), .O(N1550) );
inv1 gate( .a(N6),.O(N6_NOT) );
inv1 gate( .a(N1178),.O(N1178_NOT));
and2 gate( .a(N6_NOT), .b(p45), .O(EX111) );
and2 gate( .a(N1178_NOT), .b(EX111), .O(EX112) );
and2 gate( .a(N6), .b(p46), .O(EX113) );
and2 gate( .a(N1178_NOT), .b(EX113), .O(EX114) );
and2 gate( .a(N6_NOT), .b(p47), .O(EX115) );
and2 gate( .a(N1178), .b(EX115), .O(EX116) );
and2 gate( .a(N6), .b(p48), .O(EX117) );
and2 gate( .a(N1178), .b(EX117), .O(EX118) );
or2  gate( .a(EX112), .b(EX114), .O(EX119) );
or2  gate( .a(EX116), .b(EX119), .O(EX120) );
or2  gate( .a(EX118), .b(EX120), .O(N1551) );
and2 gate299( .a(N24), .b(N1178), .O(N1552) );
nand2 gate300( .a(N1395), .b(N1185), .O(N1553) );
nand2 gate301( .a(N1396), .b(N1397), .O(N1557) );
nand2 gate302( .a(N1398), .b(N1399), .O(N1561) );
and2 gate303( .a(N25), .b(N1200), .O(N1564) );
and2 gate304( .a(N32), .b(N1200), .O(N1565) );
and2 gate305( .a(N26), .b(N1200), .O(N1566) );
and2 gate306( .a(N33), .b(N1200), .O(N1567) );
and2 gate307( .a(N27), .b(N1205), .O(N1568) );
and2 gate308( .a(N34), .b(N1205), .O(N1569) );
and2 gate309( .a(N35), .b(N1205), .O(N1570) );
and2 gate310( .a(N28), .b(N1205), .O(N1571) );
inv1 gate311( .a(N1251), .O(N1572) );
inv1 gate312( .a(N1254), .O(N1573) );
inv1 gate313( .a(N1257), .O(N1574) );
inv1 gate314( .a(N1260), .O(N1575) );
inv1 gate315( .a(N1263), .O(N1576) );
inv1 gate316( .a(N1266), .O(N1577) );
nand2 gate317( .a(N1422), .b(N1423), .O(N1578) );
inv1 gate318( .a(N1216), .O(N1581) );
nand2 gate319( .a(N1426), .b(N1427), .O(N1582) );
inv1 gate( .a(N1424),.O(N1424_NOT) );
inv1 gate( .a(N1425),.O(N1425_NOT));
and2 gate( .a(N1424_NOT), .b(p49), .O(EX121) );
and2 gate( .a(N1425_NOT), .b(EX121), .O(EX122) );
and2 gate( .a(N1424), .b(p50), .O(EX123) );
and2 gate( .a(N1425_NOT), .b(EX123), .O(EX124) );
and2 gate( .a(N1424_NOT), .b(p51), .O(EX125) );
and2 gate( .a(N1425), .b(EX125), .O(EX126) );
and2 gate( .a(N1424), .b(p52), .O(EX127) );
and2 gate( .a(N1425), .b(EX127), .O(EX128) );
or2  gate( .a(EX122), .b(EX124), .O(EX129) );
or2  gate( .a(EX126), .b(EX129), .O(EX130) );
or2  gate( .a(EX128), .b(EX130), .O(N1585) );
nand2 gate321( .a(N1440), .b(N1441), .O(N1588) );
and2 gate322( .a(N1449), .b(N1450), .O(N1591) );
or4 gate323( .a(N1451), .b(N1452), .c(N1453), .d(N1064), .O(N1596) );
or4 gate324( .a(N1454), .b(N1455), .c(N1456), .d(N1065), .O(N1600) );
or4 gate325( .a(N1457), .b(N1458), .c(N1459), .d(N1066), .O(N1606) );
or4 gate326( .a(N1460), .b(N1461), .c(N1462), .d(N1067), .O(N1612) );
or4 gate327( .a(N1463), .b(N1464), .c(N1465), .d(N1068), .O(N1615) );
or4 gate328( .a(N1466), .b(N1467), .c(N1468), .d(N1097), .O(N1619) );
or4 gate329( .a(N1469), .b(N1470), .c(N1471), .d(N1098), .O(N1624) );
or4 gate330( .a(N1472), .b(N1473), .c(N1474), .d(N1099), .O(N1628) );
or4 gate331( .a(N1475), .b(N1476), .c(N1477), .d(N1100), .O(N1631) );
or4 gate332( .a(N1478), .b(N1479), .c(N1480), .d(N1101), .O(N1634) );
or4 gate333( .a(N1481), .b(N1482), .c(N1483), .d(N1124), .O(N1637) );
or4 gate334( .a(N1484), .b(N1485), .c(N1486), .d(N1125), .O(N1642) );
or4 gate335( .a(N1487), .b(N1488), .c(N1489), .d(N1126), .O(N1647) );
or4 gate336( .a(N1490), .b(N1491), .c(N1492), .d(N1127), .O(N1651) );
or4 gate337( .a(N1493), .b(N1494), .c(N1495), .d(N1128), .O(N1656) );
or4 gate338( .a(N1532), .b(N1533), .c(N1534), .d(N1169), .O(N1676) );
or4 gate339( .a(N1535), .b(N1536), .c(N1537), .d(N1170), .O(N1681) );
or4 gate340( .a(N1538), .b(N1539), .c(N1540), .d(N1171), .O(N1686) );
or4 gate341( .a(N1541), .b(N1542), .c(N1543), .d(N1172), .O(N1690) );
or4 gate342( .a(N1529), .b(N1530), .c(N1531), .d(N1168), .O(N1708) );
buf1 gate343( .a(N1591), .O(N1726) );
inv1 gate344( .a(N1502), .O(N1770) );
inv1 gate345( .a(N1506), .O(N1773) );
inv1 gate346( .a(N1513), .O(N1776) );
inv1 gate347( .a(N1516), .O(N1777) );
buf1 gate348( .a(N1510), .O(N1778) );
buf1 gate349( .a(N1510), .O(N1781) );
and3 gate350( .a(N1133), .b(N1129), .c(N1513), .O(N1784) );
and3 gate351( .a(N1499), .b(N1496), .c(N1516), .O(N1785) );
inv1 gate352( .a(N1553), .O(N1795) );
inv1 gate353( .a(N1557), .O(N1798) );
buf1 gate354( .a(N1561), .O(N1801) );
buf1 gate355( .a(N1561), .O(N1804) );
inv1 gate356( .a(N1588), .O(N1807) );
inv1 gate357( .a(N1578), .O(N1808) );
nand2 gate358( .a(N1578), .b(N1581), .O(N1809) );
inv1 gate359( .a(N1582), .O(N1810) );
inv1 gate360( .a(N1585), .O(N1811) );
and2 gate361( .a(N1596), .b(N241), .O(N1813) );
inv1 gate( .a(N1606),.O(N1606_NOT) );
inv1 gate( .a(N241),.O(N241_NOT));
and2 gate( .a(N1606_NOT), .b(p53), .O(EX131) );
and2 gate( .a(N241_NOT), .b(EX131), .O(EX132) );
and2 gate( .a(N1606), .b(p54), .O(EX133) );
and2 gate( .a(N241_NOT), .b(EX133), .O(EX134) );
and2 gate( .a(N1606_NOT), .b(p55), .O(EX135) );
and2 gate( .a(N241), .b(EX135), .O(EX136) );
and2 gate( .a(N1606), .b(p56), .O(EX137) );
and2 gate( .a(N241), .b(EX137), .O(EX138) );
or2  gate( .a(EX132), .b(EX134), .O(EX139) );
or2  gate( .a(EX136), .b(EX139), .O(EX140) );
or2  gate( .a(EX138), .b(EX140), .O(N1814) );
and2 gate363( .a(N1600), .b(N241), .O(N1815) );
inv1 gate364( .a(N1642), .O(N1816) );
inv1 gate365( .a(N1647), .O(N1817) );
inv1 gate366( .a(N1637), .O(N1818) );
inv1 gate367( .a(N1624), .O(N1819) );
inv1 gate368( .a(N1619), .O(N1820) );
inv1 gate369( .a(N1615), .O(N1821) );
and4 gate370( .a(N496), .b(N224), .c(N36), .d(N1591), .O(N1822) );
and4 gate371( .a(N496), .b(N224), .c(N1591), .d(N486), .O(N1823) );
buf1 gate372( .a(N1596), .O(N1824) );
inv1 gate373( .a(N1606), .O(N1827) );
and2 gate374( .a(N1600), .b(N537), .O(N1830) );
and2 gate375( .a(N1606), .b(N537), .O(N1831) );
and2 gate376( .a(N1619), .b(N246), .O(N1832) );
inv1 gate377( .a(N1596), .O(N1833) );
inv1 gate378( .a(N1600), .O(N1836) );
inv1 gate379( .a(N1606), .O(N1841) );
buf1 gate380( .a(N1612), .O(N1848) );
buf1 gate381( .a(N1615), .O(N1852) );
buf1 gate382( .a(N1619), .O(N1856) );
buf1 gate383( .a(N1624), .O(N1863) );
buf1 gate384( .a(N1628), .O(N1870) );
buf1 gate385( .a(N1631), .O(N1875) );
buf1 gate386( .a(N1634), .O(N1880) );
nand2 gate387( .a(N727), .b(N1651), .O(N1885) );
nand2 gate388( .a(N730), .b(N1656), .O(N1888) );
buf1 gate389( .a(N1686), .O(N1891) );
and2 gate390( .a(N1637), .b(N425), .O(N1894) );
inv1 gate391( .a(N1642), .O(N1897) );
and3 gate392( .a(N1496), .b(N1133), .c(N1776), .O(N1908) );
and3 gate393( .a(N1129), .b(N1499), .c(N1777), .O(N1909) );
and2 gate394( .a(N1600), .b(N637), .O(N1910) );
inv1 gate( .a(N1606),.O(N1606_NOT) );
inv1 gate( .a(N637),.O(N637_NOT));
and2 gate( .a(N1606_NOT), .b(p57), .O(EX141) );
and2 gate( .a(N637_NOT), .b(EX141), .O(EX142) );
and2 gate( .a(N1606), .b(p58), .O(EX143) );
and2 gate( .a(N637_NOT), .b(EX143), .O(EX144) );
and2 gate( .a(N1606_NOT), .b(p59), .O(EX145) );
and2 gate( .a(N637), .b(EX145), .O(EX146) );
and2 gate( .a(N1606), .b(p60), .O(EX147) );
and2 gate( .a(N637), .b(EX147), .O(EX148) );
or2  gate( .a(EX142), .b(EX144), .O(EX149) );
or2  gate( .a(EX146), .b(EX149), .O(EX150) );
or2  gate( .a(EX148), .b(EX150), .O(N1911) );
inv1 gate( .a(N1612),.O(N1612_NOT) );
inv1 gate( .a(N637),.O(N637_NOT));
and2 gate( .a(N1612_NOT), .b(p61), .O(EX151) );
and2 gate( .a(N637_NOT), .b(EX151), .O(EX152) );
and2 gate( .a(N1612), .b(p62), .O(EX153) );
and2 gate( .a(N637_NOT), .b(EX153), .O(EX154) );
and2 gate( .a(N1612_NOT), .b(p63), .O(EX155) );
and2 gate( .a(N637), .b(EX155), .O(EX156) );
and2 gate( .a(N1612), .b(p64), .O(EX157) );
and2 gate( .a(N637), .b(EX157), .O(EX158) );
or2  gate( .a(EX152), .b(EX154), .O(EX159) );
or2  gate( .a(EX156), .b(EX159), .O(EX160) );
or2  gate( .a(EX158), .b(EX160), .O(N1912) );
and2 gate397( .a(N1615), .b(N637), .O(N1913) );
inv1 gate( .a(N1619),.O(N1619_NOT) );
inv1 gate( .a(N643),.O(N643_NOT));
and2 gate( .a(N1619_NOT), .b(p65), .O(EX161) );
and2 gate( .a(N643_NOT), .b(EX161), .O(EX162) );
and2 gate( .a(N1619), .b(p66), .O(EX163) );
and2 gate( .a(N643_NOT), .b(EX163), .O(EX164) );
and2 gate( .a(N1619_NOT), .b(p67), .O(EX165) );
and2 gate( .a(N643), .b(EX165), .O(EX166) );
and2 gate( .a(N1619), .b(p68), .O(EX167) );
and2 gate( .a(N643), .b(EX167), .O(EX168) );
or2  gate( .a(EX162), .b(EX164), .O(EX169) );
or2  gate( .a(EX166), .b(EX169), .O(EX170) );
or2  gate( .a(EX168), .b(EX170), .O(N1914) );
and2 gate399( .a(N1624), .b(N643), .O(N1915) );
and2 gate400( .a(N1628), .b(N643), .O(N1916) );
inv1 gate( .a(N1631),.O(N1631_NOT) );
inv1 gate( .a(N643),.O(N643_NOT));
and2 gate( .a(N1631_NOT), .b(p69), .O(EX171) );
and2 gate( .a(N643_NOT), .b(EX171), .O(EX172) );
and2 gate( .a(N1631), .b(p70), .O(EX173) );
and2 gate( .a(N643_NOT), .b(EX173), .O(EX174) );
and2 gate( .a(N1631_NOT), .b(p71), .O(EX175) );
and2 gate( .a(N643), .b(EX175), .O(EX176) );
and2 gate( .a(N1631), .b(p72), .O(EX177) );
and2 gate( .a(N643), .b(EX177), .O(EX178) );
or2  gate( .a(EX172), .b(EX174), .O(EX179) );
or2  gate( .a(EX176), .b(EX179), .O(EX180) );
or2  gate( .a(EX178), .b(EX180), .O(N1917) );
inv1 gate( .a(N1634),.O(N1634_NOT) );
inv1 gate( .a(N643),.O(N643_NOT));
and2 gate( .a(N1634_NOT), .b(p73), .O(EX181) );
and2 gate( .a(N643_NOT), .b(EX181), .O(EX182) );
and2 gate( .a(N1634), .b(p74), .O(EX183) );
and2 gate( .a(N643_NOT), .b(EX183), .O(EX184) );
and2 gate( .a(N1634_NOT), .b(p75), .O(EX185) );
and2 gate( .a(N643), .b(EX185), .O(EX186) );
and2 gate( .a(N1634), .b(p76), .O(EX187) );
and2 gate( .a(N643), .b(EX187), .O(EX188) );
or2  gate( .a(EX182), .b(EX184), .O(EX189) );
or2  gate( .a(EX186), .b(EX189), .O(EX190) );
or2  gate( .a(EX188), .b(EX190), .O(N1918) );
inv1 gate403( .a(N1708), .O(N1919) );
inv1 gate( .a(N1676),.O(N1676_NOT) );
inv1 gate( .a(N693),.O(N693_NOT));
and2 gate( .a(N1676_NOT), .b(p77), .O(EX191) );
and2 gate( .a(N693_NOT), .b(EX191), .O(EX192) );
and2 gate( .a(N1676), .b(p78), .O(EX193) );
and2 gate( .a(N693_NOT), .b(EX193), .O(EX194) );
and2 gate( .a(N1676_NOT), .b(p79), .O(EX195) );
and2 gate( .a(N693), .b(EX195), .O(EX196) );
and2 gate( .a(N1676), .b(p80), .O(EX197) );
and2 gate( .a(N693), .b(EX197), .O(EX198) );
or2  gate( .a(EX192), .b(EX194), .O(EX199) );
or2  gate( .a(EX196), .b(EX199), .O(EX200) );
or2  gate( .a(EX198), .b(EX200), .O(N1928) );
and2 gate405( .a(N1681), .b(N693), .O(N1929) );
and2 gate406( .a(N1686), .b(N693), .O(N1930) );
and2 gate407( .a(N1690), .b(N693), .O(N1931) );
inv1 gate( .a(N1637),.O(N1637_NOT) );
inv1 gate( .a(N699),.O(N699_NOT));
and2 gate( .a(N1637_NOT), .b(p81), .O(EX201) );
and2 gate( .a(N699_NOT), .b(EX201), .O(EX202) );
and2 gate( .a(N1637), .b(p82), .O(EX203) );
and2 gate( .a(N699_NOT), .b(EX203), .O(EX204) );
and2 gate( .a(N1637_NOT), .b(p83), .O(EX205) );
and2 gate( .a(N699), .b(EX205), .O(EX206) );
and2 gate( .a(N1637), .b(p84), .O(EX207) );
and2 gate( .a(N699), .b(EX207), .O(EX208) );
or2  gate( .a(EX202), .b(EX204), .O(EX209) );
or2  gate( .a(EX206), .b(EX209), .O(EX210) );
or2  gate( .a(EX208), .b(EX210), .O(N1932) );
and2 gate409( .a(N1642), .b(N699), .O(N1933) );
inv1 gate( .a(N1647),.O(N1647_NOT) );
inv1 gate( .a(N699),.O(N699_NOT));
and2 gate( .a(N1647_NOT), .b(p85), .O(EX211) );
and2 gate( .a(N699_NOT), .b(EX211), .O(EX212) );
and2 gate( .a(N1647), .b(p86), .O(EX213) );
and2 gate( .a(N699_NOT), .b(EX213), .O(EX214) );
and2 gate( .a(N1647_NOT), .b(p87), .O(EX215) );
and2 gate( .a(N699), .b(EX215), .O(EX216) );
and2 gate( .a(N1647), .b(p88), .O(EX217) );
and2 gate( .a(N699), .b(EX217), .O(EX218) );
or2  gate( .a(EX212), .b(EX214), .O(EX219) );
or2  gate( .a(EX216), .b(EX219), .O(EX220) );
or2  gate( .a(EX218), .b(EX220), .O(N1934) );
and2 gate411( .a(N1651), .b(N699), .O(N1935) );
buf1 gate412( .a(N1600), .O(N1936) );
nand2 gate413( .a(N1216), .b(N1808), .O(N1939) );
nand2 gate414( .a(N1585), .b(N1810), .O(N1940) );
nand2 gate415( .a(N1582), .b(N1811), .O(N1941) );
buf1 gate416( .a(N1676), .O(N1942) );
buf1 gate417( .a(N1686), .O(N1945) );
buf1 gate418( .a(N1681), .O(N1948) );
buf1 gate419( .a(N1637), .O(N1951) );
buf1 gate420( .a(N1690), .O(N1954) );
buf1 gate421( .a(N1647), .O(N1957) );
buf1 gate422( .a(N1642), .O(N1960) );
buf1 gate423( .a(N1656), .O(N1963) );
buf1 gate424( .a(N1651), .O(N1966) );
inv1 gate( .a(N533),.O(N533_NOT) );
inv1 gate( .a(N1815),.O(N1815_NOT));
and2 gate( .a(N533_NOT), .b(p89), .O(EX221) );
and2 gate( .a(N1815_NOT), .b(EX221), .O(EX222) );
and2 gate( .a(N533), .b(p90), .O(EX223) );
and2 gate( .a(N1815_NOT), .b(EX223), .O(EX224) );
and2 gate( .a(N533_NOT), .b(p91), .O(EX225) );
and2 gate( .a(N1815), .b(EX225), .O(EX226) );
and2 gate( .a(N533), .b(p92), .O(EX227) );
and2 gate( .a(N1815), .b(EX227), .O(EX228) );
or2  gate( .a(EX222), .b(EX224), .O(EX229) );
or2  gate( .a(EX226), .b(EX229), .O(EX230) );
or2  gate( .a(EX228), .b(EX230), .O(N1969) );
inv1 gate426( .a(N1822), .O(N1970) );
inv1 gate427( .a(N1823), .O(N1971) );
buf1 gate428( .a(N1848), .O(N2010) );
buf1 gate429( .a(N1852), .O(N2012) );
buf1 gate430( .a(N1856), .O(N2014) );
buf1 gate431( .a(N1863), .O(N2016) );
buf1 gate432( .a(N1870), .O(N2018) );
buf1 gate433( .a(N1875), .O(N2020) );
buf1 gate434( .a(N1880), .O(N2022) );
inv1 gate435( .a(N1778), .O(N2028) );
inv1 gate436( .a(N1781), .O(N2029) );
nor2 gate437( .a(N1908), .b(N1784), .O(N2030) );
inv1 gate( .a(N1909),.O(N1909_NOT) );
inv1 gate( .a(N1785),.O(N1785_NOT));
and2 gate( .a(N1909_NOT), .b(p93), .O(EX231) );
and2 gate( .a(N1785_NOT), .b(EX231), .O(EX232) );
and2 gate( .a(N1909), .b(p94), .O(EX233) );
and2 gate( .a(N1785_NOT), .b(EX233), .O(EX234) );
and2 gate( .a(N1909_NOT), .b(p95), .O(EX235) );
and2 gate( .a(N1785), .b(EX235), .O(EX236) );
and2 gate( .a(N1909), .b(p96), .O(EX237) );
and2 gate( .a(N1785), .b(EX237), .O(EX238) );
or2  gate( .a(EX232), .b(EX234), .O(EX239) );
or2  gate( .a(EX236), .b(EX239), .O(EX240) );
or2  gate( .a(EX238), .b(EX240), .O(N2031) );
and3 gate439( .a(N1506), .b(N1502), .c(N1778), .O(N2032) );
and3 gate440( .a(N1773), .b(N1770), .c(N1781), .O(N2033) );
or2 gate441( .a(N1571), .b(N1935), .O(N2034) );
inv1 gate442( .a(N1801), .O(N2040) );
inv1 gate443( .a(N1804), .O(N2041) );
and3 gate444( .a(N1557), .b(N1553), .c(N1801), .O(N2042) );
and3 gate445( .a(N1798), .b(N1795), .c(N1804), .O(N2043) );
nand2 gate446( .a(N1939), .b(N1809), .O(N2046) );
nand2 gate447( .a(N1940), .b(N1941), .O(N2049) );
or2 gate448( .a(N1544), .b(N1910), .O(N2052) );
or2 gate449( .a(N1545), .b(N1911), .O(N2055) );
or2 gate450( .a(N1546), .b(N1912), .O(N2058) );
inv1 gate( .a(N1547),.O(N1547_NOT) );
inv1 gate( .a(N1913),.O(N1913_NOT));
and2 gate( .a(N1547_NOT), .b(p97), .O(EX241) );
and2 gate( .a(N1913_NOT), .b(EX241), .O(EX242) );
and2 gate( .a(N1547), .b(p98), .O(EX243) );
and2 gate( .a(N1913_NOT), .b(EX243), .O(EX244) );
and2 gate( .a(N1547_NOT), .b(p99), .O(EX245) );
and2 gate( .a(N1913), .b(EX245), .O(EX246) );
and2 gate( .a(N1547), .b(p100), .O(EX247) );
and2 gate( .a(N1913), .b(EX247), .O(EX248) );
or2  gate( .a(EX242), .b(EX244), .O(EX249) );
or2  gate( .a(EX246), .b(EX249), .O(EX250) );
or2  gate( .a(EX248), .b(EX250), .O(N2061) );
or2 gate452( .a(N1548), .b(N1914), .O(N2064) );
or2 gate453( .a(N1549), .b(N1915), .O(N2067) );
or2 gate454( .a(N1550), .b(N1916), .O(N2070) );
or2 gate455( .a(N1551), .b(N1917), .O(N2073) );
or2 gate456( .a(N1552), .b(N1918), .O(N2076) );
or2 gate457( .a(N1564), .b(N1928), .O(N2079) );
or2 gate458( .a(N1565), .b(N1929), .O(N2095) );
or2 gate459( .a(N1566), .b(N1930), .O(N2098) );
or2 gate460( .a(N1567), .b(N1931), .O(N2101) );
inv1 gate( .a(N1568),.O(N1568_NOT) );
inv1 gate( .a(N1932),.O(N1932_NOT));
and2 gate( .a(N1568_NOT), .b(p101), .O(EX251) );
and2 gate( .a(N1932_NOT), .b(EX251), .O(EX252) );
and2 gate( .a(N1568), .b(p102), .O(EX253) );
and2 gate( .a(N1932_NOT), .b(EX253), .O(EX254) );
and2 gate( .a(N1568_NOT), .b(p103), .O(EX255) );
and2 gate( .a(N1932), .b(EX255), .O(EX256) );
and2 gate( .a(N1568), .b(p104), .O(EX257) );
and2 gate( .a(N1932), .b(EX257), .O(EX258) );
or2  gate( .a(EX252), .b(EX254), .O(EX259) );
or2  gate( .a(EX256), .b(EX259), .O(EX260) );
or2  gate( .a(EX258), .b(EX260), .O(N2104) );
or2 gate462( .a(N1569), .b(N1933), .O(N2107) );
or2 gate463( .a(N1570), .b(N1934), .O(N2110) );
and3 gate464( .a(N1897), .b(N1894), .c(N40), .O(N2113) );
inv1 gate465( .a(N1894), .O(N2119) );
nand2 gate466( .a(N408), .b(N1827), .O(N2120) );
inv1 gate( .a(N1824),.O(N1824_NOT) );
inv1 gate( .a(N537),.O(N537_NOT));
and2 gate( .a(N1824_NOT), .b(p105), .O(EX261) );
and2 gate( .a(N537_NOT), .b(EX261), .O(EX262) );
and2 gate( .a(N1824), .b(p106), .O(EX263) );
and2 gate( .a(N537_NOT), .b(EX263), .O(EX264) );
and2 gate( .a(N1824_NOT), .b(p107), .O(EX265) );
and2 gate( .a(N537), .b(EX265), .O(EX266) );
and2 gate( .a(N1824), .b(p108), .O(EX267) );
and2 gate( .a(N537), .b(EX267), .O(EX268) );
or2  gate( .a(EX262), .b(EX264), .O(EX269) );
or2  gate( .a(EX266), .b(EX269), .O(EX270) );
or2  gate( .a(EX268), .b(EX270), .O(N2125) );
and2 gate468( .a(N1852), .b(N246), .O(N2126) );
and2 gate469( .a(N1848), .b(N537), .O(N2127) );
inv1 gate470( .a(N1848), .O(N2128) );
inv1 gate471( .a(N1852), .O(N2135) );
inv1 gate472( .a(N1863), .O(N2141) );
inv1 gate473( .a(N1870), .O(N2144) );
inv1 gate474( .a(N1875), .O(N2147) );
inv1 gate475( .a(N1880), .O(N2150) );
and2 gate476( .a(N727), .b(N1885), .O(N2153) );
and2 gate477( .a(N1885), .b(N1651), .O(N2154) );
and2 gate478( .a(N730), .b(N1888), .O(N2155) );
and2 gate479( .a(N1888), .b(N1656), .O(N2156) );
and3 gate480( .a(N1770), .b(N1506), .c(N2028), .O(N2157) );
and3 gate481( .a(N1502), .b(N1773), .c(N2029), .O(N2158) );
inv1 gate482( .a(N1942), .O(N2171) );
nand2 gate483( .a(N1942), .b(N1919), .O(N2172) );
inv1 gate484( .a(N1945), .O(N2173) );
inv1 gate485( .a(N1948), .O(N2174) );
inv1 gate486( .a(N1951), .O(N2175) );
inv1 gate487( .a(N1954), .O(N2176) );
and3 gate488( .a(N1795), .b(N1557), .c(N2040), .O(N2177) );
and3 gate489( .a(N1553), .b(N1798), .c(N2041), .O(N2178) );
buf1 gate490( .a(N1836), .O(N2185) );
buf1 gate491( .a(N1833), .O(N2188) );
buf1 gate492( .a(N1841), .O(N2191) );
inv1 gate493( .a(N1856), .O(N2194) );
inv1 gate494( .a(N1827), .O(N2197) );
inv1 gate495( .a(N1936), .O(N2200) );
buf1 gate496( .a(N1836), .O(N2201) );
buf1 gate497( .a(N1833), .O(N2204) );
buf1 gate498( .a(N1841), .O(N2207) );
buf1 gate499( .a(N1824), .O(N2210) );
buf1 gate500( .a(N1841), .O(N2213) );
buf1 gate501( .a(N1841), .O(N2216) );
nand2 gate502( .a(N2031), .b(N2030), .O(N2219) );
inv1 gate503( .a(N1957), .O(N2234) );
inv1 gate504( .a(N1960), .O(N2235) );
inv1 gate505( .a(N1963), .O(N2236) );
inv1 gate506( .a(N1966), .O(N2237) );
and3 gate507( .a(N40), .b(N1897), .c(N2119), .O(N2250) );
or2 gate508( .a(N1831), .b(N2126), .O(N2266) );
or2 gate509( .a(N2127), .b(N1832), .O(N2269) );
or2 gate510( .a(N2153), .b(N2154), .O(N2291) );
or2 gate511( .a(N2155), .b(N2156), .O(N2294) );
inv1 gate( .a(N2157),.O(N2157_NOT) );
inv1 gate( .a(N2032),.O(N2032_NOT));
and2 gate( .a(N2157_NOT), .b(p109), .O(EX271) );
and2 gate( .a(N2032_NOT), .b(EX271), .O(EX272) );
and2 gate( .a(N2157), .b(p110), .O(EX273) );
and2 gate( .a(N2032_NOT), .b(EX273), .O(EX274) );
and2 gate( .a(N2157_NOT), .b(p111), .O(EX275) );
and2 gate( .a(N2032), .b(EX275), .O(EX276) );
and2 gate( .a(N2157), .b(p112), .O(EX277) );
and2 gate( .a(N2032), .b(EX277), .O(EX278) );
or2  gate( .a(EX272), .b(EX274), .O(EX279) );
or2  gate( .a(EX276), .b(EX279), .O(EX280) );
or2  gate( .a(EX278), .b(EX280), .O(N2297) );
nor2 gate513( .a(N2158), .b(N2033), .O(N2298) );
inv1 gate514( .a(N2046), .O(N2300) );
inv1 gate515( .a(N2049), .O(N2301) );
inv1 gate( .a(N2052),.O(N2052_NOT) );
inv1 gate( .a(N1519),.O(N1519_NOT));
and2 gate( .a(N2052_NOT), .b(p113), .O(EX281) );
and2 gate( .a(N1519_NOT), .b(EX281), .O(EX282) );
and2 gate( .a(N2052), .b(p114), .O(EX283) );
and2 gate( .a(N1519_NOT), .b(EX283), .O(EX284) );
and2 gate( .a(N2052_NOT), .b(p115), .O(EX285) );
and2 gate( .a(N1519), .b(EX285), .O(EX286) );
and2 gate( .a(N2052), .b(p116), .O(EX287) );
and2 gate( .a(N1519), .b(EX287), .O(EX288) );
or2  gate( .a(EX282), .b(EX284), .O(EX289) );
or2  gate( .a(EX286), .b(EX289), .O(EX290) );
or2  gate( .a(EX288), .b(EX290), .O(N2302) );
inv1 gate517( .a(N2052), .O(N2303) );
inv1 gate( .a(N2055),.O(N2055_NOT) );
inv1 gate( .a(N1520),.O(N1520_NOT));
and2 gate( .a(N2055_NOT), .b(p117), .O(EX291) );
and2 gate( .a(N1520_NOT), .b(EX291), .O(EX292) );
and2 gate( .a(N2055), .b(p118), .O(EX293) );
and2 gate( .a(N1520_NOT), .b(EX293), .O(EX294) );
and2 gate( .a(N2055_NOT), .b(p119), .O(EX295) );
and2 gate( .a(N1520), .b(EX295), .O(EX296) );
and2 gate( .a(N2055), .b(p120), .O(EX297) );
and2 gate( .a(N1520), .b(EX297), .O(EX298) );
or2  gate( .a(EX292), .b(EX294), .O(EX299) );
or2  gate( .a(EX296), .b(EX299), .O(EX300) );
or2  gate( .a(EX298), .b(EX300), .O(N2304) );
inv1 gate519( .a(N2055), .O(N2305) );
nand2 gate520( .a(N2058), .b(N1521), .O(N2306) );
inv1 gate521( .a(N2058), .O(N2307) );
nand2 gate522( .a(N2061), .b(N1522), .O(N2308) );
inv1 gate523( .a(N2061), .O(N2309) );
nand2 gate524( .a(N2064), .b(N1523), .O(N2310) );
inv1 gate525( .a(N2064), .O(N2311) );
nand2 gate526( .a(N2067), .b(N1524), .O(N2312) );
inv1 gate527( .a(N2067), .O(N2313) );
nand2 gate528( .a(N2070), .b(N1525), .O(N2314) );
inv1 gate529( .a(N2070), .O(N2315) );
nand2 gate530( .a(N2073), .b(N1526), .O(N2316) );
inv1 gate531( .a(N2073), .O(N2317) );
inv1 gate( .a(N2076),.O(N2076_NOT) );
inv1 gate( .a(N1527),.O(N1527_NOT));
and2 gate( .a(N2076_NOT), .b(p121), .O(EX301) );
and2 gate( .a(N1527_NOT), .b(EX301), .O(EX302) );
and2 gate( .a(N2076), .b(p122), .O(EX303) );
and2 gate( .a(N1527_NOT), .b(EX303), .O(EX304) );
and2 gate( .a(N2076_NOT), .b(p123), .O(EX305) );
and2 gate( .a(N1527), .b(EX305), .O(EX306) );
and2 gate( .a(N2076), .b(p124), .O(EX307) );
and2 gate( .a(N1527), .b(EX307), .O(EX308) );
or2  gate( .a(EX302), .b(EX304), .O(EX309) );
or2  gate( .a(EX306), .b(EX309), .O(EX310) );
or2  gate( .a(EX308), .b(EX310), .O(N2318) );
inv1 gate533( .a(N2076), .O(N2319) );
nand2 gate534( .a(N2079), .b(N1528), .O(N2320) );
inv1 gate535( .a(N2079), .O(N2321) );
nand2 gate536( .a(N1708), .b(N2171), .O(N2322) );
nand2 gate537( .a(N1948), .b(N2173), .O(N2323) );
nand2 gate538( .a(N1945), .b(N2174), .O(N2324) );
nand2 gate539( .a(N1954), .b(N2175), .O(N2325) );
nand2 gate540( .a(N1951), .b(N2176), .O(N2326) );
nor2 gate541( .a(N2177), .b(N2042), .O(N2327) );
nor2 gate542( .a(N2178), .b(N2043), .O(N2328) );
nand2 gate543( .a(N2095), .b(N1572), .O(N2329) );
inv1 gate544( .a(N2095), .O(N2330) );
inv1 gate( .a(N2098),.O(N2098_NOT) );
inv1 gate( .a(N1573),.O(N1573_NOT));
and2 gate( .a(N2098_NOT), .b(p125), .O(EX311) );
and2 gate( .a(N1573_NOT), .b(EX311), .O(EX312) );
and2 gate( .a(N2098), .b(p126), .O(EX313) );
and2 gate( .a(N1573_NOT), .b(EX313), .O(EX314) );
and2 gate( .a(N2098_NOT), .b(p127), .O(EX315) );
and2 gate( .a(N1573), .b(EX315), .O(EX316) );
and2 gate( .a(N2098), .b(p128), .O(EX317) );
and2 gate( .a(N1573), .b(EX317), .O(EX318) );
or2  gate( .a(EX312), .b(EX314), .O(EX319) );
or2  gate( .a(EX316), .b(EX319), .O(EX320) );
or2  gate( .a(EX318), .b(EX320), .O(N2331) );
inv1 gate546( .a(N2098), .O(N2332) );
nand2 gate547( .a(N2101), .b(N1574), .O(N2333) );
inv1 gate548( .a(N2101), .O(N2334) );
nand2 gate549( .a(N2104), .b(N1575), .O(N2335) );
inv1 gate550( .a(N2104), .O(N2336) );
nand2 gate551( .a(N2107), .b(N1576), .O(N2337) );
inv1 gate552( .a(N2107), .O(N2338) );
inv1 gate( .a(N2110),.O(N2110_NOT) );
inv1 gate( .a(N1577),.O(N1577_NOT));
and2 gate( .a(N2110_NOT), .b(p129), .O(EX321) );
and2 gate( .a(N1577_NOT), .b(EX321), .O(EX322) );
and2 gate( .a(N2110), .b(p130), .O(EX323) );
and2 gate( .a(N1577_NOT), .b(EX323), .O(EX324) );
and2 gate( .a(N2110_NOT), .b(p131), .O(EX325) );
and2 gate( .a(N1577), .b(EX325), .O(EX326) );
and2 gate( .a(N2110), .b(p132), .O(EX327) );
and2 gate( .a(N1577), .b(EX327), .O(EX328) );
or2  gate( .a(EX322), .b(EX324), .O(EX329) );
or2  gate( .a(EX326), .b(EX329), .O(EX330) );
or2  gate( .a(EX328), .b(EX330), .O(N2339) );
inv1 gate554( .a(N2110), .O(N2340) );
nand2 gate555( .a(N1960), .b(N2234), .O(N2354) );
nand2 gate556( .a(N1957), .b(N2235), .O(N2355) );
nand2 gate557( .a(N1966), .b(N2236), .O(N2356) );
nand2 gate558( .a(N1963), .b(N2237), .O(N2357) );
inv1 gate( .a(N2120),.O(N2120_NOT) );
inv1 gate( .a(N533),.O(N533_NOT));
and2 gate( .a(N2120_NOT), .b(p133), .O(EX331) );
and2 gate( .a(N533_NOT), .b(EX331), .O(EX332) );
and2 gate( .a(N2120), .b(p134), .O(EX333) );
and2 gate( .a(N533_NOT), .b(EX333), .O(EX334) );
and2 gate( .a(N2120_NOT), .b(p135), .O(EX335) );
and2 gate( .a(N533), .b(EX335), .O(EX336) );
and2 gate( .a(N2120), .b(p136), .O(EX337) );
and2 gate( .a(N533), .b(EX337), .O(EX338) );
or2  gate( .a(EX332), .b(EX334), .O(EX339) );
or2  gate( .a(EX336), .b(EX339), .O(EX340) );
or2  gate( .a(EX338), .b(EX340), .O(N2358) );
inv1 gate560( .a(N2113), .O(N2359) );
inv1 gate561( .a(N2185), .O(N2364) );
inv1 gate562( .a(N2188), .O(N2365) );
inv1 gate563( .a(N2191), .O(N2366) );
inv1 gate564( .a(N2194), .O(N2367) );
buf1 gate565( .a(N2120), .O(N2368) );
inv1 gate566( .a(N2201), .O(N2372) );
inv1 gate567( .a(N2204), .O(N2373) );
inv1 gate568( .a(N2207), .O(N2374) );
inv1 gate569( .a(N2210), .O(N2375) );
inv1 gate570( .a(N2213), .O(N2376) );
inv1 gate571( .a(N2113), .O(N2377) );
buf1 gate572( .a(N2113), .O(N2382) );
and2 gate573( .a(N2120), .b(N246), .O(N2386) );
buf1 gate574( .a(N2266), .O(N2387) );
buf1 gate575( .a(N2266), .O(N2388) );
buf1 gate576( .a(N2269), .O(N2389) );
buf1 gate577( .a(N2269), .O(N2390) );
buf1 gate578( .a(N2113), .O(N2391) );
inv1 gate579( .a(N2113), .O(N2395) );
nand2 gate580( .a(N2219), .b(N2300), .O(N2400) );
inv1 gate581( .a(N2216), .O(N2403) );
inv1 gate582( .a(N2219), .O(N2406) );
nand2 gate583( .a(N1219), .b(N2303), .O(N2407) );
nand2 gate584( .a(N1222), .b(N2305), .O(N2408) );
nand2 gate585( .a(N1225), .b(N2307), .O(N2409) );
inv1 gate( .a(N1228),.O(N1228_NOT) );
inv1 gate( .a(N2309),.O(N2309_NOT));
and2 gate( .a(N1228_NOT), .b(p137), .O(EX341) );
and2 gate( .a(N2309_NOT), .b(EX341), .O(EX342) );
and2 gate( .a(N1228), .b(p138), .O(EX343) );
and2 gate( .a(N2309_NOT), .b(EX343), .O(EX344) );
and2 gate( .a(N1228_NOT), .b(p139), .O(EX345) );
and2 gate( .a(N2309), .b(EX345), .O(EX346) );
and2 gate( .a(N1228), .b(p140), .O(EX347) );
and2 gate( .a(N2309), .b(EX347), .O(EX348) );
or2  gate( .a(EX342), .b(EX344), .O(EX349) );
or2  gate( .a(EX346), .b(EX349), .O(EX350) );
or2  gate( .a(EX348), .b(EX350), .O(N2410) );
nand2 gate587( .a(N1231), .b(N2311), .O(N2411) );
nand2 gate588( .a(N1234), .b(N2313), .O(N2412) );
nand2 gate589( .a(N1237), .b(N2315), .O(N2413) );
inv1 gate( .a(N1240),.O(N1240_NOT) );
inv1 gate( .a(N2317),.O(N2317_NOT));
and2 gate( .a(N1240_NOT), .b(p141), .O(EX351) );
and2 gate( .a(N2317_NOT), .b(EX351), .O(EX352) );
and2 gate( .a(N1240), .b(p142), .O(EX353) );
and2 gate( .a(N2317_NOT), .b(EX353), .O(EX354) );
and2 gate( .a(N1240_NOT), .b(p143), .O(EX355) );
and2 gate( .a(N2317), .b(EX355), .O(EX356) );
and2 gate( .a(N1240), .b(p144), .O(EX357) );
and2 gate( .a(N2317), .b(EX357), .O(EX358) );
or2  gate( .a(EX352), .b(EX354), .O(EX359) );
or2  gate( .a(EX356), .b(EX359), .O(EX360) );
or2  gate( .a(EX358), .b(EX360), .O(N2414) );
nand2 gate591( .a(N1243), .b(N2319), .O(N2415) );
nand2 gate592( .a(N1246), .b(N2321), .O(N2416) );
nand2 gate593( .a(N2322), .b(N2172), .O(N2417) );
nand2 gate594( .a(N2323), .b(N2324), .O(N2421) );
nand2 gate595( .a(N2325), .b(N2326), .O(N2425) );
nand2 gate596( .a(N1251), .b(N2330), .O(N2428) );
nand2 gate597( .a(N1254), .b(N2332), .O(N2429) );
nand2 gate598( .a(N1257), .b(N2334), .O(N2430) );
nand2 gate599( .a(N1260), .b(N2336), .O(N2431) );
nand2 gate600( .a(N1263), .b(N2338), .O(N2432) );
inv1 gate( .a(N1266),.O(N1266_NOT) );
inv1 gate( .a(N2340),.O(N2340_NOT));
and2 gate( .a(N1266_NOT), .b(p145), .O(EX361) );
and2 gate( .a(N2340_NOT), .b(EX361), .O(EX362) );
and2 gate( .a(N1266), .b(p146), .O(EX363) );
and2 gate( .a(N2340_NOT), .b(EX363), .O(EX364) );
and2 gate( .a(N1266_NOT), .b(p147), .O(EX365) );
and2 gate( .a(N2340), .b(EX365), .O(EX366) );
and2 gate( .a(N1266), .b(p148), .O(EX367) );
and2 gate( .a(N2340), .b(EX367), .O(EX368) );
or2  gate( .a(EX362), .b(EX364), .O(EX369) );
or2  gate( .a(EX366), .b(EX369), .O(EX370) );
or2  gate( .a(EX368), .b(EX370), .O(N2433) );
buf1 gate602( .a(N2128), .O(N2434) );
buf1 gate603( .a(N2135), .O(N2437) );
buf1 gate604( .a(N2144), .O(N2440) );
buf1 gate605( .a(N2141), .O(N2443) );
buf1 gate606( .a(N2150), .O(N2446) );
buf1 gate607( .a(N2147), .O(N2449) );
inv1 gate608( .a(N2197), .O(N2452) );
nand2 gate609( .a(N2197), .b(N2200), .O(N2453) );
buf1 gate610( .a(N2128), .O(N2454) );
buf1 gate611( .a(N2144), .O(N2457) );
buf1 gate612( .a(N2141), .O(N2460) );
buf1 gate613( .a(N2150), .O(N2463) );
buf1 gate614( .a(N2147), .O(N2466) );
inv1 gate615( .a(N2120), .O(N2469) );
buf1 gate616( .a(N2128), .O(N2472) );
buf1 gate617( .a(N2135), .O(N2475) );
buf1 gate618( .a(N2128), .O(N2478) );
buf1 gate619( .a(N2135), .O(N2481) );
nand2 gate620( .a(N2298), .b(N2297), .O(N2484) );
nand2 gate621( .a(N2356), .b(N2357), .O(N2487) );
nand2 gate622( .a(N2354), .b(N2355), .O(N2490) );
nand2 gate623( .a(N2328), .b(N2327), .O(N2493) );
or2 gate624( .a(N2358), .b(N1814), .O(N2496) );
nand2 gate625( .a(N2188), .b(N2364), .O(N2503) );
nand2 gate626( .a(N2185), .b(N2365), .O(N2504) );
nand2 gate627( .a(N2204), .b(N2372), .O(N2510) );
nand2 gate628( .a(N2201), .b(N2373), .O(N2511) );
or2 gate629( .a(N1830), .b(N2386), .O(N2521) );
nand2 gate630( .a(N2046), .b(N2406), .O(N2528) );
inv1 gate631( .a(N2291), .O(N2531) );
inv1 gate632( .a(N2294), .O(N2534) );
buf1 gate633( .a(N2250), .O(N2537) );
buf1 gate634( .a(N2250), .O(N2540) );
inv1 gate( .a(N2302),.O(N2302_NOT) );
inv1 gate( .a(N2407),.O(N2407_NOT));
and2 gate( .a(N2302_NOT), .b(p149), .O(EX371) );
and2 gate( .a(N2407_NOT), .b(EX371), .O(EX372) );
and2 gate( .a(N2302), .b(p150), .O(EX373) );
and2 gate( .a(N2407_NOT), .b(EX373), .O(EX374) );
and2 gate( .a(N2302_NOT), .b(p151), .O(EX375) );
and2 gate( .a(N2407), .b(EX375), .O(EX376) );
and2 gate( .a(N2302), .b(p152), .O(EX377) );
and2 gate( .a(N2407), .b(EX377), .O(EX378) );
or2  gate( .a(EX372), .b(EX374), .O(EX379) );
or2  gate( .a(EX376), .b(EX379), .O(EX380) );
or2  gate( .a(EX378), .b(EX380), .O(N2544) );
nand2 gate636( .a(N2304), .b(N2408), .O(N2545) );
nand2 gate637( .a(N2306), .b(N2409), .O(N2546) );
inv1 gate( .a(N2308),.O(N2308_NOT) );
inv1 gate( .a(N2410),.O(N2410_NOT));
and2 gate( .a(N2308_NOT), .b(p153), .O(EX381) );
and2 gate( .a(N2410_NOT), .b(EX381), .O(EX382) );
and2 gate( .a(N2308), .b(p154), .O(EX383) );
and2 gate( .a(N2410_NOT), .b(EX383), .O(EX384) );
and2 gate( .a(N2308_NOT), .b(p155), .O(EX385) );
and2 gate( .a(N2410), .b(EX385), .O(EX386) );
and2 gate( .a(N2308), .b(p156), .O(EX387) );
and2 gate( .a(N2410), .b(EX387), .O(EX388) );
or2  gate( .a(EX382), .b(EX384), .O(EX389) );
or2  gate( .a(EX386), .b(EX389), .O(EX390) );
or2  gate( .a(EX388), .b(EX390), .O(N2547) );
inv1 gate( .a(N2310),.O(N2310_NOT) );
inv1 gate( .a(N2411),.O(N2411_NOT));
and2 gate( .a(N2310_NOT), .b(p157), .O(EX391) );
and2 gate( .a(N2411_NOT), .b(EX391), .O(EX392) );
and2 gate( .a(N2310), .b(p158), .O(EX393) );
and2 gate( .a(N2411_NOT), .b(EX393), .O(EX394) );
and2 gate( .a(N2310_NOT), .b(p159), .O(EX395) );
and2 gate( .a(N2411), .b(EX395), .O(EX396) );
and2 gate( .a(N2310), .b(p160), .O(EX397) );
and2 gate( .a(N2411), .b(EX397), .O(EX398) );
or2  gate( .a(EX392), .b(EX394), .O(EX399) );
or2  gate( .a(EX396), .b(EX399), .O(EX400) );
or2  gate( .a(EX398), .b(EX400), .O(N2548) );
nand2 gate640( .a(N2312), .b(N2412), .O(N2549) );
nand2 gate641( .a(N2314), .b(N2413), .O(N2550) );
nand2 gate642( .a(N2316), .b(N2414), .O(N2551) );
inv1 gate( .a(N2318),.O(N2318_NOT) );
inv1 gate( .a(N2415),.O(N2415_NOT));
and2 gate( .a(N2318_NOT), .b(p161), .O(EX401) );
and2 gate( .a(N2415_NOT), .b(EX401), .O(EX402) );
and2 gate( .a(N2318), .b(p162), .O(EX403) );
and2 gate( .a(N2415_NOT), .b(EX403), .O(EX404) );
and2 gate( .a(N2318_NOT), .b(p163), .O(EX405) );
and2 gate( .a(N2415), .b(EX405), .O(EX406) );
and2 gate( .a(N2318), .b(p164), .O(EX407) );
and2 gate( .a(N2415), .b(EX407), .O(EX408) );
or2  gate( .a(EX402), .b(EX404), .O(EX409) );
or2  gate( .a(EX406), .b(EX409), .O(EX410) );
or2  gate( .a(EX408), .b(EX410), .O(N2552) );
nand2 gate644( .a(N2320), .b(N2416), .O(N2553) );
nand2 gate645( .a(N2329), .b(N2428), .O(N2563) );
nand2 gate646( .a(N2331), .b(N2429), .O(N2564) );
nand2 gate647( .a(N2333), .b(N2430), .O(N2565) );
nand2 gate648( .a(N2335), .b(N2431), .O(N2566) );
nand2 gate649( .a(N2337), .b(N2432), .O(N2567) );
nand2 gate650( .a(N2339), .b(N2433), .O(N2568) );
inv1 gate( .a(N1936),.O(N1936_NOT) );
inv1 gate( .a(N2452),.O(N2452_NOT));
and2 gate( .a(N1936_NOT), .b(p165), .O(EX411) );
and2 gate( .a(N2452_NOT), .b(EX411), .O(EX412) );
and2 gate( .a(N1936), .b(p166), .O(EX413) );
and2 gate( .a(N2452_NOT), .b(EX413), .O(EX414) );
and2 gate( .a(N1936_NOT), .b(p167), .O(EX415) );
and2 gate( .a(N2452), .b(EX415), .O(EX416) );
and2 gate( .a(N1936), .b(p168), .O(EX417) );
and2 gate( .a(N2452), .b(EX417), .O(EX418) );
or2  gate( .a(EX412), .b(EX414), .O(EX419) );
or2  gate( .a(EX416), .b(EX419), .O(EX420) );
or2  gate( .a(EX418), .b(EX420), .O(N2579) );
buf1 gate652( .a(N2359), .O(N2603) );
and2 gate653( .a(N1880), .b(N2377), .O(N2607) );
inv1 gate( .a(N1676),.O(N1676_NOT) );
inv1 gate( .a(N2377),.O(N2377_NOT));
and2 gate( .a(N1676_NOT), .b(p169), .O(EX421) );
and2 gate( .a(N2377_NOT), .b(EX421), .O(EX422) );
and2 gate( .a(N1676), .b(p170), .O(EX423) );
and2 gate( .a(N2377_NOT), .b(EX423), .O(EX424) );
and2 gate( .a(N1676_NOT), .b(p171), .O(EX425) );
and2 gate( .a(N2377), .b(EX425), .O(EX426) );
and2 gate( .a(N1676), .b(p172), .O(EX427) );
and2 gate( .a(N2377), .b(EX427), .O(EX428) );
or2  gate( .a(EX422), .b(EX424), .O(EX429) );
or2  gate( .a(EX426), .b(EX429), .O(EX430) );
or2  gate( .a(EX428), .b(EX430), .O(N2608) );
inv1 gate( .a(N1681),.O(N1681_NOT) );
inv1 gate( .a(N2377),.O(N2377_NOT));
and2 gate( .a(N1681_NOT), .b(p173), .O(EX431) );
and2 gate( .a(N2377_NOT), .b(EX431), .O(EX432) );
and2 gate( .a(N1681), .b(p174), .O(EX433) );
and2 gate( .a(N2377_NOT), .b(EX433), .O(EX434) );
and2 gate( .a(N1681_NOT), .b(p175), .O(EX435) );
and2 gate( .a(N2377), .b(EX435), .O(EX436) );
and2 gate( .a(N1681), .b(p176), .O(EX437) );
and2 gate( .a(N2377), .b(EX437), .O(EX438) );
or2  gate( .a(EX432), .b(EX434), .O(EX439) );
or2  gate( .a(EX436), .b(EX439), .O(EX440) );
or2  gate( .a(EX438), .b(EX440), .O(N2609) );
and2 gate656( .a(N1891), .b(N2377), .O(N2610) );
and2 gate657( .a(N1856), .b(N2382), .O(N2611) );
and2 gate658( .a(N1863), .b(N2382), .O(N2612) );
nand2 gate659( .a(N2503), .b(N2504), .O(N2613) );
inv1 gate660( .a(N2434), .O(N2617) );
nand2 gate661( .a(N2434), .b(N2366), .O(N2618) );
nand2 gate662( .a(N2437), .b(N2367), .O(N2619) );
inv1 gate663( .a(N2437), .O(N2620) );
inv1 gate664( .a(N2368), .O(N2621) );
nand2 gate665( .a(N2510), .b(N2511), .O(N2624) );
inv1 gate666( .a(N2454), .O(N2628) );
nand2 gate667( .a(N2454), .b(N2374), .O(N2629) );
inv1 gate668( .a(N2472), .O(N2630) );
and2 gate669( .a(N1856), .b(N2391), .O(N2631) );
inv1 gate( .a(N1863),.O(N1863_NOT) );
inv1 gate( .a(N2391),.O(N2391_NOT));
and2 gate( .a(N1863_NOT), .b(p177), .O(EX441) );
and2 gate( .a(N2391_NOT), .b(EX441), .O(EX442) );
and2 gate( .a(N1863), .b(p178), .O(EX443) );
and2 gate( .a(N2391_NOT), .b(EX443), .O(EX444) );
and2 gate( .a(N1863_NOT), .b(p179), .O(EX445) );
and2 gate( .a(N2391), .b(EX445), .O(EX446) );
and2 gate( .a(N1863), .b(p180), .O(EX447) );
and2 gate( .a(N2391), .b(EX447), .O(EX448) );
or2  gate( .a(EX442), .b(EX444), .O(EX449) );
or2  gate( .a(EX446), .b(EX449), .O(EX450) );
or2  gate( .a(EX448), .b(EX450), .O(N2632) );
inv1 gate( .a(N1880),.O(N1880_NOT) );
inv1 gate( .a(N2395),.O(N2395_NOT));
and2 gate( .a(N1880_NOT), .b(p181), .O(EX451) );
and2 gate( .a(N2395_NOT), .b(EX451), .O(EX452) );
and2 gate( .a(N1880), .b(p182), .O(EX453) );
and2 gate( .a(N2395_NOT), .b(EX453), .O(EX454) );
and2 gate( .a(N1880_NOT), .b(p183), .O(EX455) );
and2 gate( .a(N2395), .b(EX455), .O(EX456) );
and2 gate( .a(N1880), .b(p184), .O(EX457) );
and2 gate( .a(N2395), .b(EX457), .O(EX458) );
or2  gate( .a(EX452), .b(EX454), .O(EX459) );
or2  gate( .a(EX456), .b(EX459), .O(EX460) );
or2  gate( .a(EX458), .b(EX460), .O(N2633) );
and2 gate672( .a(N1676), .b(N2395), .O(N2634) );
and2 gate673( .a(N1681), .b(N2395), .O(N2635) );
and2 gate674( .a(N1891), .b(N2395), .O(N2636) );
inv1 gate675( .a(N2382), .O(N2638) );
buf1 gate676( .a(N2521), .O(N2643) );
buf1 gate677( .a(N2521), .O(N2644) );
inv1 gate678( .a(N2475), .O(N2645) );
inv1 gate679( .a(N2391), .O(N2646) );
nand2 gate680( .a(N2528), .b(N2400), .O(N2652) );
inv1 gate681( .a(N2478), .O(N2655) );
inv1 gate682( .a(N2481), .O(N2656) );
buf1 gate683( .a(N2359), .O(N2659) );
inv1 gate684( .a(N2484), .O(N2663) );
nand2 gate685( .a(N2484), .b(N2301), .O(N2664) );
inv1 gate686( .a(N2553), .O(N2665) );
inv1 gate687( .a(N2552), .O(N2666) );
inv1 gate688( .a(N2551), .O(N2667) );
inv1 gate689( .a(N2550), .O(N2668) );
inv1 gate690( .a(N2549), .O(N2669) );
inv1 gate691( .a(N2548), .O(N2670) );
inv1 gate692( .a(N2547), .O(N2671) );
inv1 gate693( .a(N2546), .O(N2672) );
inv1 gate694( .a(N2545), .O(N2673) );
inv1 gate695( .a(N2544), .O(N2674) );
inv1 gate696( .a(N2568), .O(N2675) );
inv1 gate697( .a(N2567), .O(N2676) );
inv1 gate698( .a(N2566), .O(N2677) );
inv1 gate699( .a(N2565), .O(N2678) );
inv1 gate700( .a(N2564), .O(N2679) );
inv1 gate701( .a(N2563), .O(N2680) );
inv1 gate702( .a(N2417), .O(N2681) );
inv1 gate703( .a(N2421), .O(N2684) );
buf1 gate704( .a(N2425), .O(N2687) );
buf1 gate705( .a(N2425), .O(N2690) );
inv1 gate706( .a(N2493), .O(N2693) );
nand2 gate707( .a(N2493), .b(N1807), .O(N2694) );
inv1 gate708( .a(N2440), .O(N2695) );
inv1 gate709( .a(N2443), .O(N2696) );
inv1 gate710( .a(N2446), .O(N2697) );
inv1 gate711( .a(N2449), .O(N2698) );
inv1 gate712( .a(N2457), .O(N2699) );
inv1 gate713( .a(N2460), .O(N2700) );
inv1 gate714( .a(N2463), .O(N2701) );
inv1 gate715( .a(N2466), .O(N2702) );
nand2 gate716( .a(N2579), .b(N2453), .O(N2703) );
inv1 gate717( .a(N2469), .O(N2706) );
inv1 gate718( .a(N2487), .O(N2707) );
inv1 gate719( .a(N2490), .O(N2708) );
inv1 gate( .a(N2294),.O(N2294_NOT) );
inv1 gate( .a(N2534),.O(N2534_NOT));
and2 gate( .a(N2294_NOT), .b(p185), .O(EX461) );
and2 gate( .a(N2534_NOT), .b(EX461), .O(EX462) );
and2 gate( .a(N2294), .b(p186), .O(EX463) );
and2 gate( .a(N2534_NOT), .b(EX463), .O(EX464) );
and2 gate( .a(N2294_NOT), .b(p187), .O(EX465) );
and2 gate( .a(N2534), .b(EX465), .O(EX466) );
and2 gate( .a(N2294), .b(p188), .O(EX467) );
and2 gate( .a(N2534), .b(EX467), .O(EX468) );
or2  gate( .a(EX462), .b(EX464), .O(EX469) );
or2  gate( .a(EX466), .b(EX469), .O(EX470) );
or2  gate( .a(EX468), .b(EX470), .O(N2709) );
and2 gate721( .a(N2291), .b(N2531), .O(N2710) );
nand2 gate722( .a(N2191), .b(N2617), .O(N2719) );
nand2 gate723( .a(N2194), .b(N2620), .O(N2720) );
nand2 gate724( .a(N2207), .b(N2628), .O(N2726) );
buf1 gate725( .a(N2537), .O(N2729) );
buf1 gate726( .a(N2537), .O(N2738) );
inv1 gate727( .a(N2652), .O(N2743) );
nand2 gate728( .a(N2049), .b(N2663), .O(N2747) );
and5 gate729( .a(N2665), .b(N2666), .c(N2667), .d(N2668), .e(N2669), .O(N2748) );
and5 gate730( .a(N2670), .b(N2671), .c(N2672), .d(N2673), .e(N2674), .O(N2749) );
and2 gate731( .a(N2034), .b(N2675), .O(N2750) );
and5 gate732( .a(N2676), .b(N2677), .c(N2678), .d(N2679), .e(N2680), .O(N2751) );
nand2 gate733( .a(N1588), .b(N2693), .O(N2760) );
buf1 gate734( .a(N2540), .O(N2761) );
buf1 gate735( .a(N2540), .O(N2766) );
inv1 gate( .a(N2443),.O(N2443_NOT) );
inv1 gate( .a(N2695),.O(N2695_NOT));
and2 gate( .a(N2443_NOT), .b(p189), .O(EX471) );
and2 gate( .a(N2695_NOT), .b(EX471), .O(EX472) );
and2 gate( .a(N2443), .b(p190), .O(EX473) );
and2 gate( .a(N2695_NOT), .b(EX473), .O(EX474) );
and2 gate( .a(N2443_NOT), .b(p191), .O(EX475) );
and2 gate( .a(N2695), .b(EX475), .O(EX476) );
and2 gate( .a(N2443), .b(p192), .O(EX477) );
and2 gate( .a(N2695), .b(EX477), .O(EX478) );
or2  gate( .a(EX472), .b(EX474), .O(EX479) );
or2  gate( .a(EX476), .b(EX479), .O(EX480) );
or2  gate( .a(EX478), .b(EX480), .O(N2771) );
nand2 gate737( .a(N2440), .b(N2696), .O(N2772) );
nand2 gate738( .a(N2449), .b(N2697), .O(N2773) );
nand2 gate739( .a(N2446), .b(N2698), .O(N2774) );
nand2 gate740( .a(N2460), .b(N2699), .O(N2775) );
nand2 gate741( .a(N2457), .b(N2700), .O(N2776) );
nand2 gate742( .a(N2466), .b(N2701), .O(N2777) );
nand2 gate743( .a(N2463), .b(N2702), .O(N2778) );
nand2 gate744( .a(N2490), .b(N2707), .O(N2781) );
nand2 gate745( .a(N2487), .b(N2708), .O(N2782) );
inv1 gate( .a(N2709),.O(N2709_NOT) );
inv1 gate( .a(N2534),.O(N2534_NOT));
and2 gate( .a(N2709_NOT), .b(p193), .O(EX481) );
and2 gate( .a(N2534_NOT), .b(EX481), .O(EX482) );
and2 gate( .a(N2709), .b(p194), .O(EX483) );
and2 gate( .a(N2534_NOT), .b(EX483), .O(EX484) );
and2 gate( .a(N2709_NOT), .b(p195), .O(EX485) );
and2 gate( .a(N2534), .b(EX485), .O(EX486) );
and2 gate( .a(N2709), .b(p196), .O(EX487) );
and2 gate( .a(N2534), .b(EX487), .O(EX488) );
or2  gate( .a(EX482), .b(EX484), .O(EX489) );
or2  gate( .a(EX486), .b(EX489), .O(EX490) );
or2  gate( .a(EX488), .b(EX490), .O(N2783) );
or2 gate747( .a(N2710), .b(N2531), .O(N2784) );
inv1 gate( .a(N1856),.O(N1856_NOT) );
inv1 gate( .a(N2638),.O(N2638_NOT));
and2 gate( .a(N1856_NOT), .b(p197), .O(EX491) );
and2 gate( .a(N2638_NOT), .b(EX491), .O(EX492) );
and2 gate( .a(N1856), .b(p198), .O(EX493) );
and2 gate( .a(N2638_NOT), .b(EX493), .O(EX494) );
and2 gate( .a(N1856_NOT), .b(p199), .O(EX495) );
and2 gate( .a(N2638), .b(EX495), .O(EX496) );
and2 gate( .a(N1856), .b(p200), .O(EX497) );
and2 gate( .a(N2638), .b(EX497), .O(EX498) );
or2  gate( .a(EX492), .b(EX494), .O(EX499) );
or2  gate( .a(EX496), .b(EX499), .O(EX500) );
or2  gate( .a(EX498), .b(EX500), .O(N2789) );
and2 gate749( .a(N1863), .b(N2638), .O(N2790) );
and2 gate750( .a(N1870), .b(N2638), .O(N2791) );
and2 gate751( .a(N1875), .b(N2638), .O(N2792) );
inv1 gate752( .a(N2613), .O(N2793) );
nand2 gate753( .a(N2719), .b(N2618), .O(N2796) );
nand2 gate754( .a(N2619), .b(N2720), .O(N2800) );
inv1 gate755( .a(N2624), .O(N2803) );
nand2 gate756( .a(N2726), .b(N2629), .O(N2806) );
and2 gate757( .a(N1856), .b(N2646), .O(N2809) );
and2 gate758( .a(N1863), .b(N2646), .O(N2810) );
and2 gate759( .a(N1870), .b(N2646), .O(N2811) );
and2 gate760( .a(N1875), .b(N2646), .O(N2812) );
and2 gate761( .a(N2743), .b(N14), .O(N2817) );
buf1 gate762( .a(N2603), .O(N2820) );
nand2 gate763( .a(N2747), .b(N2664), .O(N2826) );
and2 gate764( .a(N2748), .b(N2749), .O(N2829) );
inv1 gate( .a(N2750),.O(N2750_NOT) );
inv1 gate( .a(N2751),.O(N2751_NOT));
and2 gate( .a(N2750_NOT), .b(p201), .O(EX501) );
and2 gate( .a(N2751_NOT), .b(EX501), .O(EX502) );
and2 gate( .a(N2750), .b(p202), .O(EX503) );
and2 gate( .a(N2751_NOT), .b(EX503), .O(EX504) );
and2 gate( .a(N2750_NOT), .b(p203), .O(EX505) );
and2 gate( .a(N2751), .b(EX505), .O(EX506) );
and2 gate( .a(N2750), .b(p204), .O(EX507) );
and2 gate( .a(N2751), .b(EX507), .O(EX508) );
or2  gate( .a(EX502), .b(EX504), .O(EX509) );
or2  gate( .a(EX506), .b(EX509), .O(EX510) );
or2  gate( .a(EX508), .b(EX510), .O(N2830) );
buf1 gate766( .a(N2659), .O(N2831) );
inv1 gate767( .a(N2687), .O(N2837) );
inv1 gate768( .a(N2690), .O(N2838) );
and3 gate769( .a(N2421), .b(N2417), .c(N2687), .O(N2839) );
and3 gate770( .a(N2684), .b(N2681), .c(N2690), .O(N2840) );
nand2 gate771( .a(N2760), .b(N2694), .O(N2841) );
buf1 gate772( .a(N2603), .O(N2844) );
buf1 gate773( .a(N2603), .O(N2854) );
buf1 gate774( .a(N2659), .O(N2859) );
buf1 gate775( .a(N2659), .O(N2869) );
nand2 gate776( .a(N2773), .b(N2774), .O(N2874) );
nand2 gate777( .a(N2771), .b(N2772), .O(N2877) );
inv1 gate778( .a(N2703), .O(N2880) );
nand2 gate779( .a(N2703), .b(N2706), .O(N2881) );
nand2 gate780( .a(N2777), .b(N2778), .O(N2882) );
nand2 gate781( .a(N2775), .b(N2776), .O(N2885) );
nand2 gate782( .a(N2781), .b(N2782), .O(N2888) );
nand2 gate783( .a(N2783), .b(N2784), .O(N2891) );
and2 gate784( .a(N2607), .b(N2729), .O(N2894) );
and2 gate785( .a(N2608), .b(N2729), .O(N2895) );
and2 gate786( .a(N2609), .b(N2729), .O(N2896) );
and2 gate787( .a(N2610), .b(N2729), .O(N2897) );
or2 gate788( .a(N2789), .b(N2611), .O(N2898) );
or2 gate789( .a(N2790), .b(N2612), .O(N2899) );
and2 gate790( .a(N2791), .b(N1037), .O(N2900) );
and2 gate791( .a(N2792), .b(N1037), .O(N2901) );
or2 gate792( .a(N2809), .b(N2631), .O(N2914) );
or2 gate793( .a(N2810), .b(N2632), .O(N2915) );
inv1 gate( .a(N2811),.O(N2811_NOT) );
inv1 gate( .a(N1070),.O(N1070_NOT));
and2 gate( .a(N2811_NOT), .b(p205), .O(EX511) );
and2 gate( .a(N1070_NOT), .b(EX511), .O(EX512) );
and2 gate( .a(N2811), .b(p206), .O(EX513) );
and2 gate( .a(N1070_NOT), .b(EX513), .O(EX514) );
and2 gate( .a(N2811_NOT), .b(p207), .O(EX515) );
and2 gate( .a(N1070), .b(EX515), .O(EX516) );
and2 gate( .a(N2811), .b(p208), .O(EX517) );
and2 gate( .a(N1070), .b(EX517), .O(EX518) );
or2  gate( .a(EX512), .b(EX514), .O(EX519) );
or2  gate( .a(EX516), .b(EX519), .O(EX520) );
or2  gate( .a(EX518), .b(EX520), .O(N2916) );
and2 gate795( .a(N2812), .b(N1070), .O(N2917) );
and2 gate796( .a(N2633), .b(N2738), .O(N2918) );
and2 gate797( .a(N2634), .b(N2738), .O(N2919) );
and2 gate798( .a(N2635), .b(N2738), .O(N2920) );
inv1 gate( .a(N2636),.O(N2636_NOT) );
inv1 gate( .a(N2738),.O(N2738_NOT));
and2 gate( .a(N2636_NOT), .b(p209), .O(EX521) );
and2 gate( .a(N2738_NOT), .b(EX521), .O(EX522) );
and2 gate( .a(N2636), .b(p210), .O(EX523) );
and2 gate( .a(N2738_NOT), .b(EX523), .O(EX524) );
and2 gate( .a(N2636_NOT), .b(p211), .O(EX525) );
and2 gate( .a(N2738), .b(EX525), .O(EX526) );
and2 gate( .a(N2636), .b(p212), .O(EX527) );
and2 gate( .a(N2738), .b(EX527), .O(EX528) );
or2  gate( .a(EX522), .b(EX524), .O(EX529) );
or2  gate( .a(EX526), .b(EX529), .O(EX530) );
or2  gate( .a(EX528), .b(EX530), .O(N2921) );
buf1 gate800( .a(N2817), .O(N2925) );
and3 gate801( .a(N2829), .b(N2830), .c(N1302), .O(N2931) );
and3 gate802( .a(N2681), .b(N2421), .c(N2837), .O(N2938) );
and3 gate803( .a(N2417), .b(N2684), .c(N2838), .O(N2939) );
nand2 gate804( .a(N2469), .b(N2880), .O(N2963) );
inv1 gate805( .a(N2841), .O(N2970) );
inv1 gate806( .a(N2826), .O(N2971) );
inv1 gate807( .a(N2894), .O(N2972) );
inv1 gate808( .a(N2895), .O(N2975) );
inv1 gate809( .a(N2896), .O(N2978) );
inv1 gate810( .a(N2897), .O(N2981) );
and2 gate811( .a(N2898), .b(N1037), .O(N2984) );
and2 gate812( .a(N2899), .b(N1037), .O(N2985) );
inv1 gate813( .a(N2900), .O(N2986) );
inv1 gate814( .a(N2901), .O(N2989) );
inv1 gate815( .a(N2796), .O(N2992) );
buf1 gate816( .a(N2800), .O(N2995) );
buf1 gate817( .a(N2800), .O(N2998) );
buf1 gate818( .a(N2806), .O(N3001) );
buf1 gate819( .a(N2806), .O(N3004) );
and2 gate820( .a(N574), .b(N2820), .O(N3007) );
and2 gate821( .a(N2914), .b(N1070), .O(N3008) );
and2 gate822( .a(N2915), .b(N1070), .O(N3009) );
inv1 gate823( .a(N2916), .O(N3010) );
inv1 gate824( .a(N2917), .O(N3013) );
inv1 gate825( .a(N2918), .O(N3016) );
inv1 gate826( .a(N2919), .O(N3019) );
inv1 gate827( .a(N2920), .O(N3022) );
inv1 gate828( .a(N2921), .O(N3025) );
inv1 gate829( .a(N2817), .O(N3028) );
and2 gate830( .a(N574), .b(N2831), .O(N3029) );
inv1 gate831( .a(N2820), .O(N3030) );
and2 gate832( .a(N578), .b(N2820), .O(N3035) );
and2 gate833( .a(N655), .b(N2820), .O(N3036) );
and2 gate834( .a(N659), .b(N2820), .O(N3037) );
buf1 gate835( .a(N2931), .O(N3038) );
inv1 gate836( .a(N2831), .O(N3039) );
inv1 gate( .a(N578),.O(N578_NOT) );
inv1 gate( .a(N2831),.O(N2831_NOT));
and2 gate( .a(N578_NOT), .b(p213), .O(EX531) );
and2 gate( .a(N2831_NOT), .b(EX531), .O(EX532) );
and2 gate( .a(N578), .b(p214), .O(EX533) );
and2 gate( .a(N2831_NOT), .b(EX533), .O(EX534) );
and2 gate( .a(N578_NOT), .b(p215), .O(EX535) );
and2 gate( .a(N2831), .b(EX535), .O(EX536) );
and2 gate( .a(N578), .b(p216), .O(EX537) );
and2 gate( .a(N2831), .b(EX537), .O(EX538) );
or2  gate( .a(EX532), .b(EX534), .O(EX539) );
or2  gate( .a(EX536), .b(EX539), .O(EX540) );
or2  gate( .a(EX538), .b(EX540), .O(N3044) );
and2 gate838( .a(N655), .b(N2831), .O(N3045) );
and2 gate839( .a(N659), .b(N2831), .O(N3046) );
inv1 gate( .a(N2938),.O(N2938_NOT) );
inv1 gate( .a(N2839),.O(N2839_NOT));
and2 gate( .a(N2938_NOT), .b(p217), .O(EX541) );
and2 gate( .a(N2839_NOT), .b(EX541), .O(EX542) );
and2 gate( .a(N2938), .b(p218), .O(EX543) );
and2 gate( .a(N2839_NOT), .b(EX543), .O(EX544) );
and2 gate( .a(N2938_NOT), .b(p219), .O(EX545) );
and2 gate( .a(N2839), .b(EX545), .O(EX546) );
and2 gate( .a(N2938), .b(p220), .O(EX547) );
and2 gate( .a(N2839), .b(EX547), .O(EX548) );
or2  gate( .a(EX542), .b(EX544), .O(EX549) );
or2  gate( .a(EX546), .b(EX549), .O(EX550) );
or2  gate( .a(EX548), .b(EX550), .O(N3047) );
nor2 gate841( .a(N2939), .b(N2840), .O(N3048) );
inv1 gate842( .a(N2888), .O(N3049) );
inv1 gate843( .a(N2844), .O(N3050) );
and2 gate844( .a(N663), .b(N2844), .O(N3053) );
and2 gate845( .a(N667), .b(N2844), .O(N3054) );
and2 gate846( .a(N671), .b(N2844), .O(N3055) );
and2 gate847( .a(N675), .b(N2844), .O(N3056) );
and2 gate848( .a(N679), .b(N2854), .O(N3057) );
and2 gate849( .a(N683), .b(N2854), .O(N3058) );
inv1 gate( .a(N687),.O(N687_NOT) );
inv1 gate( .a(N2854),.O(N2854_NOT));
and2 gate( .a(N687_NOT), .b(p221), .O(EX551) );
and2 gate( .a(N2854_NOT), .b(EX551), .O(EX552) );
and2 gate( .a(N687), .b(p222), .O(EX553) );
and2 gate( .a(N2854_NOT), .b(EX553), .O(EX554) );
and2 gate( .a(N687_NOT), .b(p223), .O(EX555) );
and2 gate( .a(N2854), .b(EX555), .O(EX556) );
and2 gate( .a(N687), .b(p224), .O(EX557) );
and2 gate( .a(N2854), .b(EX557), .O(EX558) );
or2  gate( .a(EX552), .b(EX554), .O(EX559) );
or2  gate( .a(EX556), .b(EX559), .O(EX560) );
or2  gate( .a(EX558), .b(EX560), .O(N3059) );
and2 gate851( .a(N705), .b(N2854), .O(N3060) );
inv1 gate852( .a(N2859), .O(N3061) );
inv1 gate( .a(N663),.O(N663_NOT) );
inv1 gate( .a(N2859),.O(N2859_NOT));
and2 gate( .a(N663_NOT), .b(p225), .O(EX561) );
and2 gate( .a(N2859_NOT), .b(EX561), .O(EX562) );
and2 gate( .a(N663), .b(p226), .O(EX563) );
and2 gate( .a(N2859_NOT), .b(EX563), .O(EX564) );
and2 gate( .a(N663_NOT), .b(p227), .O(EX565) );
and2 gate( .a(N2859), .b(EX565), .O(EX566) );
and2 gate( .a(N663), .b(p228), .O(EX567) );
and2 gate( .a(N2859), .b(EX567), .O(EX568) );
or2  gate( .a(EX562), .b(EX564), .O(EX569) );
or2  gate( .a(EX566), .b(EX569), .O(EX570) );
or2  gate( .a(EX568), .b(EX570), .O(N3064) );
inv1 gate( .a(N667),.O(N667_NOT) );
inv1 gate( .a(N2859),.O(N2859_NOT));
and2 gate( .a(N667_NOT), .b(p229), .O(EX571) );
and2 gate( .a(N2859_NOT), .b(EX571), .O(EX572) );
and2 gate( .a(N667), .b(p230), .O(EX573) );
and2 gate( .a(N2859_NOT), .b(EX573), .O(EX574) );
and2 gate( .a(N667_NOT), .b(p231), .O(EX575) );
and2 gate( .a(N2859), .b(EX575), .O(EX576) );
and2 gate( .a(N667), .b(p232), .O(EX577) );
and2 gate( .a(N2859), .b(EX577), .O(EX578) );
or2  gate( .a(EX572), .b(EX574), .O(EX579) );
or2  gate( .a(EX576), .b(EX579), .O(EX580) );
or2  gate( .a(EX578), .b(EX580), .O(N3065) );
and2 gate855( .a(N671), .b(N2859), .O(N3066) );
and2 gate856( .a(N675), .b(N2859), .O(N3067) );
inv1 gate( .a(N679),.O(N679_NOT) );
inv1 gate( .a(N2869),.O(N2869_NOT));
and2 gate( .a(N679_NOT), .b(p233), .O(EX581) );
and2 gate( .a(N2869_NOT), .b(EX581), .O(EX582) );
and2 gate( .a(N679), .b(p234), .O(EX583) );
and2 gate( .a(N2869_NOT), .b(EX583), .O(EX584) );
and2 gate( .a(N679_NOT), .b(p235), .O(EX585) );
and2 gate( .a(N2869), .b(EX585), .O(EX586) );
and2 gate( .a(N679), .b(p236), .O(EX587) );
and2 gate( .a(N2869), .b(EX587), .O(EX588) );
or2  gate( .a(EX582), .b(EX584), .O(EX589) );
or2  gate( .a(EX586), .b(EX589), .O(EX590) );
or2  gate( .a(EX588), .b(EX590), .O(N3068) );
and2 gate858( .a(N683), .b(N2869), .O(N3069) );
and2 gate859( .a(N687), .b(N2869), .O(N3070) );
and2 gate860( .a(N705), .b(N2869), .O(N3071) );
inv1 gate861( .a(N2874), .O(N3072) );
inv1 gate862( .a(N2877), .O(N3073) );
inv1 gate863( .a(N2882), .O(N3074) );
inv1 gate864( .a(N2885), .O(N3075) );
nand2 gate865( .a(N2881), .b(N2963), .O(N3076) );
inv1 gate866( .a(N2931), .O(N3079) );
inv1 gate867( .a(N2984), .O(N3088) );
inv1 gate868( .a(N2985), .O(N3091) );
inv1 gate869( .a(N3008), .O(N3110) );
inv1 gate870( .a(N3009), .O(N3113) );
and2 gate871( .a(N3055), .b(N1190), .O(N3137) );
inv1 gate( .a(N3056),.O(N3056_NOT) );
inv1 gate( .a(N1190),.O(N1190_NOT));
and2 gate( .a(N3056_NOT), .b(p237), .O(EX591) );
and2 gate( .a(N1190_NOT), .b(EX591), .O(EX592) );
and2 gate( .a(N3056), .b(p238), .O(EX593) );
and2 gate( .a(N1190_NOT), .b(EX593), .O(EX594) );
and2 gate( .a(N3056_NOT), .b(p239), .O(EX595) );
and2 gate( .a(N1190), .b(EX595), .O(EX596) );
and2 gate( .a(N3056), .b(p240), .O(EX597) );
and2 gate( .a(N1190), .b(EX597), .O(EX598) );
or2  gate( .a(EX592), .b(EX594), .O(EX599) );
or2  gate( .a(EX596), .b(EX599), .O(EX600) );
or2  gate( .a(EX598), .b(EX600), .O(N3140) );
and2 gate873( .a(N3057), .b(N2761), .O(N3143) );
and2 gate874( .a(N3058), .b(N2761), .O(N3146) );
inv1 gate( .a(N3059),.O(N3059_NOT) );
inv1 gate( .a(N2761),.O(N2761_NOT));
and2 gate( .a(N3059_NOT), .b(p241), .O(EX601) );
and2 gate( .a(N2761_NOT), .b(EX601), .O(EX602) );
and2 gate( .a(N3059), .b(p242), .O(EX603) );
and2 gate( .a(N2761_NOT), .b(EX603), .O(EX604) );
and2 gate( .a(N3059_NOT), .b(p243), .O(EX605) );
and2 gate( .a(N2761), .b(EX605), .O(EX606) );
and2 gate( .a(N3059), .b(p244), .O(EX607) );
and2 gate( .a(N2761), .b(EX607), .O(EX608) );
or2  gate( .a(EX602), .b(EX604), .O(EX609) );
or2  gate( .a(EX606), .b(EX609), .O(EX610) );
or2  gate( .a(EX608), .b(EX610), .O(N3149) );
and2 gate876( .a(N3060), .b(N2761), .O(N3152) );
inv1 gate( .a(N3066),.O(N3066_NOT) );
inv1 gate( .a(N1195),.O(N1195_NOT));
and2 gate( .a(N3066_NOT), .b(p245), .O(EX611) );
and2 gate( .a(N1195_NOT), .b(EX611), .O(EX612) );
and2 gate( .a(N3066), .b(p246), .O(EX613) );
and2 gate( .a(N1195_NOT), .b(EX613), .O(EX614) );
and2 gate( .a(N3066_NOT), .b(p247), .O(EX615) );
and2 gate( .a(N1195), .b(EX615), .O(EX616) );
and2 gate( .a(N3066), .b(p248), .O(EX617) );
and2 gate( .a(N1195), .b(EX617), .O(EX618) );
or2  gate( .a(EX612), .b(EX614), .O(EX619) );
or2  gate( .a(EX616), .b(EX619), .O(EX620) );
or2  gate( .a(EX618), .b(EX620), .O(N3157) );
and2 gate878( .a(N3067), .b(N1195), .O(N3160) );
and2 gate879( .a(N3068), .b(N2766), .O(N3163) );
and2 gate880( .a(N3069), .b(N2766), .O(N3166) );
and2 gate881( .a(N3070), .b(N2766), .O(N3169) );
and2 gate882( .a(N3071), .b(N2766), .O(N3172) );
nand2 gate883( .a(N2877), .b(N3072), .O(N3175) );
nand2 gate884( .a(N2874), .b(N3073), .O(N3176) );
nand2 gate885( .a(N2885), .b(N3074), .O(N3177) );
nand2 gate886( .a(N2882), .b(N3075), .O(N3178) );
nand2 gate887( .a(N3048), .b(N3047), .O(N3180) );
inv1 gate888( .a(N2995), .O(N3187) );
inv1 gate889( .a(N2998), .O(N3188) );
inv1 gate890( .a(N3001), .O(N3189) );
inv1 gate891( .a(N3004), .O(N3190) );
and3 gate892( .a(N2796), .b(N2613), .c(N2995), .O(N3191) );
and3 gate893( .a(N2992), .b(N2793), .c(N2998), .O(N3192) );
and3 gate894( .a(N2624), .b(N2368), .c(N3001), .O(N3193) );
and3 gate895( .a(N2803), .b(N2621), .c(N3004), .O(N3194) );
nand2 gate896( .a(N3076), .b(N2375), .O(N3195) );
inv1 gate897( .a(N3076), .O(N3196) );
and2 gate898( .a(N687), .b(N3030), .O(N3197) );
and2 gate899( .a(N687), .b(N3039), .O(N3208) );
inv1 gate( .a(N705),.O(N705_NOT) );
inv1 gate( .a(N3030),.O(N3030_NOT));
and2 gate( .a(N705_NOT), .b(p249), .O(EX621) );
and2 gate( .a(N3030_NOT), .b(EX621), .O(EX622) );
and2 gate( .a(N705), .b(p250), .O(EX623) );
and2 gate( .a(N3030_NOT), .b(EX623), .O(EX624) );
and2 gate( .a(N705_NOT), .b(p251), .O(EX625) );
and2 gate( .a(N3030), .b(EX625), .O(EX626) );
and2 gate( .a(N705), .b(p252), .O(EX627) );
and2 gate( .a(N3030), .b(EX627), .O(EX628) );
or2  gate( .a(EX622), .b(EX624), .O(EX629) );
or2  gate( .a(EX626), .b(EX629), .O(EX630) );
or2  gate( .a(EX628), .b(EX630), .O(N3215) );
and2 gate901( .a(N711), .b(N3030), .O(N3216) );
and2 gate902( .a(N715), .b(N3030), .O(N3217) );
and2 gate903( .a(N705), .b(N3039), .O(N3218) );
and2 gate904( .a(N711), .b(N3039), .O(N3219) );
and2 gate905( .a(N715), .b(N3039), .O(N3220) );
inv1 gate( .a(N719),.O(N719_NOT) );
inv1 gate( .a(N3050),.O(N3050_NOT));
and2 gate( .a(N719_NOT), .b(p253), .O(EX631) );
and2 gate( .a(N3050_NOT), .b(EX631), .O(EX632) );
and2 gate( .a(N719), .b(p254), .O(EX633) );
and2 gate( .a(N3050_NOT), .b(EX633), .O(EX634) );
and2 gate( .a(N719_NOT), .b(p255), .O(EX635) );
and2 gate( .a(N3050), .b(EX635), .O(EX636) );
and2 gate( .a(N719), .b(p256), .O(EX637) );
and2 gate( .a(N3050), .b(EX637), .O(EX638) );
or2  gate( .a(EX632), .b(EX634), .O(EX639) );
or2  gate( .a(EX636), .b(EX639), .O(EX640) );
or2  gate( .a(EX638), .b(EX640), .O(N3222) );
inv1 gate( .a(N723),.O(N723_NOT) );
inv1 gate( .a(N3050),.O(N3050_NOT));
and2 gate( .a(N723_NOT), .b(p257), .O(EX641) );
and2 gate( .a(N3050_NOT), .b(EX641), .O(EX642) );
and2 gate( .a(N723), .b(p258), .O(EX643) );
and2 gate( .a(N3050_NOT), .b(EX643), .O(EX644) );
and2 gate( .a(N723_NOT), .b(p259), .O(EX645) );
and2 gate( .a(N3050), .b(EX645), .O(EX646) );
and2 gate( .a(N723), .b(p260), .O(EX647) );
and2 gate( .a(N3050), .b(EX647), .O(EX648) );
or2  gate( .a(EX642), .b(EX644), .O(EX649) );
or2  gate( .a(EX646), .b(EX649), .O(EX650) );
or2  gate( .a(EX648), .b(EX650), .O(N3223) );
inv1 gate( .a(N719),.O(N719_NOT) );
inv1 gate( .a(N3061),.O(N3061_NOT));
and2 gate( .a(N719_NOT), .b(p261), .O(EX651) );
and2 gate( .a(N3061_NOT), .b(EX651), .O(EX652) );
and2 gate( .a(N719), .b(p262), .O(EX653) );
and2 gate( .a(N3061_NOT), .b(EX653), .O(EX654) );
and2 gate( .a(N719_NOT), .b(p263), .O(EX655) );
and2 gate( .a(N3061), .b(EX655), .O(EX656) );
and2 gate( .a(N719), .b(p264), .O(EX657) );
and2 gate( .a(N3061), .b(EX657), .O(EX658) );
or2  gate( .a(EX652), .b(EX654), .O(EX659) );
or2  gate( .a(EX656), .b(EX659), .O(EX660) );
or2  gate( .a(EX658), .b(EX660), .O(N3230) );
inv1 gate( .a(N723),.O(N723_NOT) );
inv1 gate( .a(N3061),.O(N3061_NOT));
and2 gate( .a(N723_NOT), .b(p265), .O(EX661) );
and2 gate( .a(N3061_NOT), .b(EX661), .O(EX662) );
and2 gate( .a(N723), .b(p266), .O(EX663) );
and2 gate( .a(N3061_NOT), .b(EX663), .O(EX664) );
and2 gate( .a(N723_NOT), .b(p267), .O(EX665) );
and2 gate( .a(N3061), .b(EX665), .O(EX666) );
and2 gate( .a(N723), .b(p268), .O(EX667) );
and2 gate( .a(N3061), .b(EX667), .O(EX668) );
or2  gate( .a(EX662), .b(EX664), .O(EX669) );
or2  gate( .a(EX666), .b(EX669), .O(EX670) );
or2  gate( .a(EX668), .b(EX670), .O(N3231) );
nand2 gate910( .a(N3175), .b(N3176), .O(N3238) );
nand2 gate911( .a(N3177), .b(N3178), .O(N3241) );
buf1 gate912( .a(N2981), .O(N3244) );
buf1 gate913( .a(N2978), .O(N3247) );
buf1 gate914( .a(N2975), .O(N3250) );
buf1 gate915( .a(N2972), .O(N3253) );
buf1 gate916( .a(N2989), .O(N3256) );
buf1 gate917( .a(N2986), .O(N3259) );
buf1 gate918( .a(N3025), .O(N3262) );
buf1 gate919( .a(N3022), .O(N3265) );
buf1 gate920( .a(N3019), .O(N3268) );
buf1 gate921( .a(N3016), .O(N3271) );
buf1 gate922( .a(N3013), .O(N3274) );
buf1 gate923( .a(N3010), .O(N3277) );
and3 gate924( .a(N2793), .b(N2796), .c(N3187), .O(N3281) );
and3 gate925( .a(N2613), .b(N2992), .c(N3188), .O(N3282) );
and3 gate926( .a(N2621), .b(N2624), .c(N3189), .O(N3283) );
and3 gate927( .a(N2368), .b(N2803), .c(N3190), .O(N3284) );
inv1 gate( .a(N2210),.O(N2210_NOT) );
inv1 gate( .a(N3196),.O(N3196_NOT));
and2 gate( .a(N2210_NOT), .b(p269), .O(EX671) );
and2 gate( .a(N3196_NOT), .b(EX671), .O(EX672) );
and2 gate( .a(N2210), .b(p270), .O(EX673) );
and2 gate( .a(N3196_NOT), .b(EX673), .O(EX674) );
and2 gate( .a(N2210_NOT), .b(p271), .O(EX675) );
and2 gate( .a(N3196), .b(EX675), .O(EX676) );
and2 gate( .a(N2210), .b(p272), .O(EX677) );
and2 gate( .a(N3196), .b(EX677), .O(EX678) );
or2  gate( .a(EX672), .b(EX674), .O(EX679) );
or2  gate( .a(EX676), .b(EX679), .O(EX680) );
or2  gate( .a(EX678), .b(EX680), .O(N3286) );
or2 gate929( .a(N3197), .b(N3007), .O(N3288) );
nand2 gate930( .a(N3180), .b(N3049), .O(N3289) );
inv1 gate( .a(N3152),.O(N3152_NOT) );
inv1 gate( .a(N2981),.O(N2981_NOT));
and2 gate( .a(N3152_NOT), .b(p273), .O(EX681) );
and2 gate( .a(N2981_NOT), .b(EX681), .O(EX682) );
and2 gate( .a(N3152), .b(p274), .O(EX683) );
and2 gate( .a(N2981_NOT), .b(EX683), .O(EX684) );
and2 gate( .a(N3152_NOT), .b(p275), .O(EX685) );
and2 gate( .a(N2981), .b(EX685), .O(EX686) );
and2 gate( .a(N3152), .b(p276), .O(EX687) );
and2 gate( .a(N2981), .b(EX687), .O(EX688) );
or2  gate( .a(EX682), .b(EX684), .O(EX689) );
or2  gate( .a(EX686), .b(EX689), .O(EX690) );
or2  gate( .a(EX688), .b(EX690), .O(N3291) );
inv1 gate( .a(N3149),.O(N3149_NOT) );
inv1 gate( .a(N2978),.O(N2978_NOT));
and2 gate( .a(N3149_NOT), .b(p277), .O(EX691) );
and2 gate( .a(N2978_NOT), .b(EX691), .O(EX692) );
and2 gate( .a(N3149), .b(p278), .O(EX693) );
and2 gate( .a(N2978_NOT), .b(EX693), .O(EX694) );
and2 gate( .a(N3149_NOT), .b(p279), .O(EX695) );
and2 gate( .a(N2978), .b(EX695), .O(EX696) );
and2 gate( .a(N3149), .b(p280), .O(EX697) );
and2 gate( .a(N2978), .b(EX697), .O(EX698) );
or2  gate( .a(EX692), .b(EX694), .O(EX699) );
or2  gate( .a(EX696), .b(EX699), .O(EX700) );
or2  gate( .a(EX698), .b(EX700), .O(N3293) );
and2 gate933( .a(N3146), .b(N2975), .O(N3295) );
and2 gate934( .a(N2972), .b(N3143), .O(N3296) );
and2 gate935( .a(N3140), .b(N2989), .O(N3299) );
and2 gate936( .a(N3137), .b(N2986), .O(N3301) );
or2 gate937( .a(N3208), .b(N3029), .O(N3302) );
inv1 gate( .a(N3172),.O(N3172_NOT) );
inv1 gate( .a(N3025),.O(N3025_NOT));
and2 gate( .a(N3172_NOT), .b(p281), .O(EX701) );
and2 gate( .a(N3025_NOT), .b(EX701), .O(EX702) );
and2 gate( .a(N3172), .b(p282), .O(EX703) );
and2 gate( .a(N3025_NOT), .b(EX703), .O(EX704) );
and2 gate( .a(N3172_NOT), .b(p283), .O(EX705) );
and2 gate( .a(N3025), .b(EX705), .O(EX706) );
and2 gate( .a(N3172), .b(p284), .O(EX707) );
and2 gate( .a(N3025), .b(EX707), .O(EX708) );
or2  gate( .a(EX702), .b(EX704), .O(EX709) );
or2  gate( .a(EX706), .b(EX709), .O(EX710) );
or2  gate( .a(EX708), .b(EX710), .O(N3304) );
and2 gate939( .a(N3169), .b(N3022), .O(N3306) );
and2 gate940( .a(N3166), .b(N3019), .O(N3308) );
and2 gate941( .a(N3016), .b(N3163), .O(N3309) );
and2 gate942( .a(N3160), .b(N3013), .O(N3312) );
and2 gate943( .a(N3157), .b(N3010), .O(N3314) );
or2 gate944( .a(N3215), .b(N3035), .O(N3315) );
or2 gate945( .a(N3216), .b(N3036), .O(N3318) );
or2 gate946( .a(N3217), .b(N3037), .O(N3321) );
or2 gate947( .a(N3218), .b(N3044), .O(N3324) );
inv1 gate( .a(N3219),.O(N3219_NOT) );
inv1 gate( .a(N3045),.O(N3045_NOT));
and2 gate( .a(N3219_NOT), .b(p285), .O(EX711) );
and2 gate( .a(N3045_NOT), .b(EX711), .O(EX712) );
and2 gate( .a(N3219), .b(p286), .O(EX713) );
and2 gate( .a(N3045_NOT), .b(EX713), .O(EX714) );
and2 gate( .a(N3219_NOT), .b(p287), .O(EX715) );
and2 gate( .a(N3045), .b(EX715), .O(EX716) );
and2 gate( .a(N3219), .b(p288), .O(EX717) );
and2 gate( .a(N3045), .b(EX717), .O(EX718) );
or2  gate( .a(EX712), .b(EX714), .O(EX719) );
or2  gate( .a(EX716), .b(EX719), .O(EX720) );
or2  gate( .a(EX718), .b(EX720), .O(N3327) );
or2 gate949( .a(N3220), .b(N3046), .O(N3330) );
inv1 gate950( .a(N3180), .O(N3333) );
or2 gate951( .a(N3222), .b(N3053), .O(N3334) );
or2 gate952( .a(N3223), .b(N3054), .O(N3335) );
or2 gate953( .a(N3230), .b(N3064), .O(N3336) );
or2 gate954( .a(N3231), .b(N3065), .O(N3337) );
buf1 gate955( .a(N3152), .O(N3340) );
buf1 gate956( .a(N3149), .O(N3344) );
buf1 gate957( .a(N3146), .O(N3348) );
buf1 gate958( .a(N3143), .O(N3352) );
buf1 gate959( .a(N3140), .O(N3356) );
buf1 gate960( .a(N3137), .O(N3360) );
buf1 gate961( .a(N3091), .O(N3364) );
buf1 gate962( .a(N3088), .O(N3367) );
buf1 gate963( .a(N3172), .O(N3370) );
buf1 gate964( .a(N3169), .O(N3374) );
buf1 gate965( .a(N3166), .O(N3378) );
buf1 gate966( .a(N3163), .O(N3382) );
buf1 gate967( .a(N3160), .O(N3386) );
buf1 gate968( .a(N3157), .O(N3390) );
buf1 gate969( .a(N3113), .O(N3394) );
buf1 gate970( .a(N3110), .O(N3397) );
inv1 gate( .a(N3195),.O(N3195_NOT) );
inv1 gate( .a(N3286),.O(N3286_NOT));
and2 gate( .a(N3195_NOT), .b(p289), .O(EX721) );
and2 gate( .a(N3286_NOT), .b(EX721), .O(EX722) );
and2 gate( .a(N3195), .b(p290), .O(EX723) );
and2 gate( .a(N3286_NOT), .b(EX723), .O(EX724) );
and2 gate( .a(N3195_NOT), .b(p291), .O(EX725) );
and2 gate( .a(N3286), .b(EX725), .O(EX726) );
and2 gate( .a(N3195), .b(p292), .O(EX727) );
and2 gate( .a(N3286), .b(EX727), .O(EX728) );
or2  gate( .a(EX722), .b(EX724), .O(EX729) );
or2  gate( .a(EX726), .b(EX729), .O(EX730) );
or2  gate( .a(EX728), .b(EX730), .O(N3400) );
nor2 gate972( .a(N3281), .b(N3191), .O(N3401) );
nor2 gate973( .a(N3282), .b(N3192), .O(N3402) );
inv1 gate( .a(N3283),.O(N3283_NOT) );
inv1 gate( .a(N3193),.O(N3193_NOT));
and2 gate( .a(N3283_NOT), .b(p293), .O(EX731) );
and2 gate( .a(N3193_NOT), .b(EX731), .O(EX732) );
and2 gate( .a(N3283), .b(p294), .O(EX733) );
and2 gate( .a(N3193_NOT), .b(EX733), .O(EX734) );
and2 gate( .a(N3283_NOT), .b(p295), .O(EX735) );
and2 gate( .a(N3193), .b(EX735), .O(EX736) );
and2 gate( .a(N3283), .b(p296), .O(EX737) );
and2 gate( .a(N3193), .b(EX737), .O(EX738) );
or2  gate( .a(EX732), .b(EX734), .O(EX739) );
or2  gate( .a(EX736), .b(EX739), .O(EX740) );
or2  gate( .a(EX738), .b(EX740), .O(N3403) );
nor2 gate975( .a(N3284), .b(N3194), .O(N3404) );
inv1 gate976( .a(N3238), .O(N3405) );
inv1 gate977( .a(N3241), .O(N3406) );
and2 gate978( .a(N3288), .b(N1836), .O(N3409) );
nand2 gate979( .a(N2888), .b(N3333), .O(N3410) );
inv1 gate980( .a(N3244), .O(N3412) );
inv1 gate981( .a(N3247), .O(N3414) );
inv1 gate982( .a(N3250), .O(N3416) );
inv1 gate983( .a(N3253), .O(N3418) );
inv1 gate984( .a(N3256), .O(N3420) );
inv1 gate985( .a(N3259), .O(N3422) );
and2 gate986( .a(N3302), .b(N1836), .O(N3428) );
inv1 gate987( .a(N3262), .O(N3430) );
inv1 gate988( .a(N3265), .O(N3432) );
inv1 gate989( .a(N3268), .O(N3434) );
inv1 gate990( .a(N3271), .O(N3436) );
inv1 gate991( .a(N3274), .O(N3438) );
inv1 gate992( .a(N3277), .O(N3440) );
and2 gate993( .a(N3334), .b(N1190), .O(N3450) );
inv1 gate( .a(N3335),.O(N3335_NOT) );
inv1 gate( .a(N1190),.O(N1190_NOT));
and2 gate( .a(N3335_NOT), .b(p297), .O(EX741) );
and2 gate( .a(N1190_NOT), .b(EX741), .O(EX742) );
and2 gate( .a(N3335), .b(p298), .O(EX743) );
and2 gate( .a(N1190_NOT), .b(EX743), .O(EX744) );
and2 gate( .a(N3335_NOT), .b(p299), .O(EX745) );
and2 gate( .a(N1190), .b(EX745), .O(EX746) );
and2 gate( .a(N3335), .b(p300), .O(EX747) );
and2 gate( .a(N1190), .b(EX747), .O(EX748) );
or2  gate( .a(EX742), .b(EX744), .O(EX749) );
or2  gate( .a(EX746), .b(EX749), .O(EX750) );
or2  gate( .a(EX748), .b(EX750), .O(N3453) );
and2 gate995( .a(N3336), .b(N1195), .O(N3456) );
and2 gate996( .a(N3337), .b(N1195), .O(N3459) );
inv1 gate( .a(N3400),.O(N3400_NOT) );
inv1 gate( .a(N533),.O(N533_NOT));
and2 gate( .a(N3400_NOT), .b(p301), .O(EX751) );
and2 gate( .a(N533_NOT), .b(EX751), .O(EX752) );
and2 gate( .a(N3400), .b(p302), .O(EX753) );
and2 gate( .a(N533_NOT), .b(EX753), .O(EX754) );
and2 gate( .a(N3400_NOT), .b(p303), .O(EX755) );
and2 gate( .a(N533), .b(EX755), .O(EX756) );
and2 gate( .a(N3400), .b(p304), .O(EX757) );
and2 gate( .a(N533), .b(EX757), .O(EX758) );
or2  gate( .a(EX752), .b(EX754), .O(EX759) );
or2  gate( .a(EX756), .b(EX759), .O(EX760) );
or2  gate( .a(EX758), .b(EX760), .O(N3478) );
and2 gate998( .a(N3318), .b(N2128), .O(N3479) );
inv1 gate( .a(N3315),.O(N3315_NOT) );
inv1 gate( .a(N1841),.O(N1841_NOT));
and2 gate( .a(N3315_NOT), .b(p305), .O(EX761) );
and2 gate( .a(N1841_NOT), .b(EX761), .O(EX762) );
and2 gate( .a(N3315), .b(p306), .O(EX763) );
and2 gate( .a(N1841_NOT), .b(EX763), .O(EX764) );
and2 gate( .a(N3315_NOT), .b(p307), .O(EX765) );
and2 gate( .a(N1841), .b(EX765), .O(EX766) );
and2 gate( .a(N3315), .b(p308), .O(EX767) );
and2 gate( .a(N1841), .b(EX767), .O(EX768) );
or2  gate( .a(EX762), .b(EX764), .O(EX769) );
or2  gate( .a(EX766), .b(EX769), .O(EX770) );
or2  gate( .a(EX768), .b(EX770), .O(N3480) );
nand2 gate1000( .a(N3410), .b(N3289), .O(N3481) );
inv1 gate1001( .a(N3340), .O(N3482) );
nand2 gate1002( .a(N3340), .b(N3412), .O(N3483) );
inv1 gate1003( .a(N3344), .O(N3484) );
inv1 gate( .a(N3344),.O(N3344_NOT) );
inv1 gate( .a(N3414),.O(N3414_NOT));
and2 gate( .a(N3344_NOT), .b(p309), .O(EX771) );
and2 gate( .a(N3414_NOT), .b(EX771), .O(EX772) );
and2 gate( .a(N3344), .b(p310), .O(EX773) );
and2 gate( .a(N3414_NOT), .b(EX773), .O(EX774) );
and2 gate( .a(N3344_NOT), .b(p311), .O(EX775) );
and2 gate( .a(N3414), .b(EX775), .O(EX776) );
and2 gate( .a(N3344), .b(p312), .O(EX777) );
and2 gate( .a(N3414), .b(EX777), .O(EX778) );
or2  gate( .a(EX772), .b(EX774), .O(EX779) );
or2  gate( .a(EX776), .b(EX779), .O(EX780) );
or2  gate( .a(EX778), .b(EX780), .O(N3485) );
inv1 gate1005( .a(N3348), .O(N3486) );
nand2 gate1006( .a(N3348), .b(N3416), .O(N3487) );
inv1 gate1007( .a(N3352), .O(N3488) );
nand2 gate1008( .a(N3352), .b(N3418), .O(N3489) );
inv1 gate1009( .a(N3356), .O(N3490) );
nand2 gate1010( .a(N3356), .b(N3420), .O(N3491) );
inv1 gate1011( .a(N3360), .O(N3492) );
nand2 gate1012( .a(N3360), .b(N3422), .O(N3493) );
inv1 gate1013( .a(N3364), .O(N3494) );
inv1 gate1014( .a(N3367), .O(N3496) );
and2 gate1015( .a(N3321), .b(N2135), .O(N3498) );
and2 gate1016( .a(N3327), .b(N2128), .O(N3499) );
and2 gate1017( .a(N3324), .b(N1841), .O(N3500) );
inv1 gate1018( .a(N3370), .O(N3501) );
inv1 gate( .a(N3370),.O(N3370_NOT) );
inv1 gate( .a(N3430),.O(N3430_NOT));
and2 gate( .a(N3370_NOT), .b(p313), .O(EX781) );
and2 gate( .a(N3430_NOT), .b(EX781), .O(EX782) );
and2 gate( .a(N3370), .b(p314), .O(EX783) );
and2 gate( .a(N3430_NOT), .b(EX783), .O(EX784) );
and2 gate( .a(N3370_NOT), .b(p315), .O(EX785) );
and2 gate( .a(N3430), .b(EX785), .O(EX786) );
and2 gate( .a(N3370), .b(p316), .O(EX787) );
and2 gate( .a(N3430), .b(EX787), .O(EX788) );
or2  gate( .a(EX782), .b(EX784), .O(EX789) );
or2  gate( .a(EX786), .b(EX789), .O(EX790) );
or2  gate( .a(EX788), .b(EX790), .O(N3502) );
inv1 gate1020( .a(N3374), .O(N3503) );
nand2 gate1021( .a(N3374), .b(N3432), .O(N3504) );
inv1 gate1022( .a(N3378), .O(N3505) );
inv1 gate( .a(N3378),.O(N3378_NOT) );
inv1 gate( .a(N3434),.O(N3434_NOT));
and2 gate( .a(N3378_NOT), .b(p317), .O(EX791) );
and2 gate( .a(N3434_NOT), .b(EX791), .O(EX792) );
and2 gate( .a(N3378), .b(p318), .O(EX793) );
and2 gate( .a(N3434_NOT), .b(EX793), .O(EX794) );
and2 gate( .a(N3378_NOT), .b(p319), .O(EX795) );
and2 gate( .a(N3434), .b(EX795), .O(EX796) );
and2 gate( .a(N3378), .b(p320), .O(EX797) );
and2 gate( .a(N3434), .b(EX797), .O(EX798) );
or2  gate( .a(EX792), .b(EX794), .O(EX799) );
or2  gate( .a(EX796), .b(EX799), .O(EX800) );
or2  gate( .a(EX798), .b(EX800), .O(N3506) );
inv1 gate1024( .a(N3382), .O(N3507) );
nand2 gate1025( .a(N3382), .b(N3436), .O(N3508) );
inv1 gate1026( .a(N3386), .O(N3509) );
nand2 gate1027( .a(N3386), .b(N3438), .O(N3510) );
inv1 gate1028( .a(N3390), .O(N3511) );
nand2 gate1029( .a(N3390), .b(N3440), .O(N3512) );
inv1 gate1030( .a(N3394), .O(N3513) );
inv1 gate1031( .a(N3397), .O(N3515) );
and2 gate1032( .a(N3330), .b(N2135), .O(N3517) );
nand2 gate1033( .a(N3402), .b(N3401), .O(N3522) );
inv1 gate( .a(N3404),.O(N3404_NOT) );
inv1 gate( .a(N3403),.O(N3403_NOT));
and2 gate( .a(N3404_NOT), .b(p321), .O(EX801) );
and2 gate( .a(N3403_NOT), .b(EX801), .O(EX802) );
and2 gate( .a(N3404), .b(p322), .O(EX803) );
and2 gate( .a(N3403_NOT), .b(EX803), .O(EX804) );
and2 gate( .a(N3404_NOT), .b(p323), .O(EX805) );
and2 gate( .a(N3403), .b(EX805), .O(EX806) );
and2 gate( .a(N3404), .b(p324), .O(EX807) );
and2 gate( .a(N3403), .b(EX807), .O(EX808) );
or2  gate( .a(EX802), .b(EX804), .O(EX809) );
or2  gate( .a(EX806), .b(EX809), .O(EX810) );
or2  gate( .a(EX808), .b(EX810), .O(N3525) );
buf1 gate1035( .a(N3318), .O(N3528) );
buf1 gate1036( .a(N3315), .O(N3531) );
buf1 gate1037( .a(N3321), .O(N3534) );
buf1 gate1038( .a(N3327), .O(N3537) );
buf1 gate1039( .a(N3324), .O(N3540) );
buf1 gate1040( .a(N3330), .O(N3543) );
or2 gate1041( .a(N3478), .b(N1813), .O(N3546) );
inv1 gate1042( .a(N3481), .O(N3551) );
nand2 gate1043( .a(N3244), .b(N3482), .O(N3552) );
nand2 gate1044( .a(N3247), .b(N3484), .O(N3553) );
inv1 gate( .a(N3250),.O(N3250_NOT) );
inv1 gate( .a(N3486),.O(N3486_NOT));
and2 gate( .a(N3250_NOT), .b(p325), .O(EX811) );
and2 gate( .a(N3486_NOT), .b(EX811), .O(EX812) );
and2 gate( .a(N3250), .b(p326), .O(EX813) );
and2 gate( .a(N3486_NOT), .b(EX813), .O(EX814) );
and2 gate( .a(N3250_NOT), .b(p327), .O(EX815) );
and2 gate( .a(N3486), .b(EX815), .O(EX816) );
and2 gate( .a(N3250), .b(p328), .O(EX817) );
and2 gate( .a(N3486), .b(EX817), .O(EX818) );
or2  gate( .a(EX812), .b(EX814), .O(EX819) );
or2  gate( .a(EX816), .b(EX819), .O(EX820) );
or2  gate( .a(EX818), .b(EX820), .O(N3554) );
nand2 gate1046( .a(N3253), .b(N3488), .O(N3555) );
nand2 gate1047( .a(N3256), .b(N3490), .O(N3556) );
nand2 gate1048( .a(N3259), .b(N3492), .O(N3557) );
and2 gate1049( .a(N3453), .b(N3091), .O(N3558) );
and2 gate1050( .a(N3450), .b(N3088), .O(N3559) );
nand2 gate1051( .a(N3262), .b(N3501), .O(N3563) );
nand2 gate1052( .a(N3265), .b(N3503), .O(N3564) );
nand2 gate1053( .a(N3268), .b(N3505), .O(N3565) );
nand2 gate1054( .a(N3271), .b(N3507), .O(N3566) );
nand2 gate1055( .a(N3274), .b(N3509), .O(N3567) );
nand2 gate1056( .a(N3277), .b(N3511), .O(N3568) );
and2 gate1057( .a(N3459), .b(N3113), .O(N3569) );
and2 gate1058( .a(N3456), .b(N3110), .O(N3570) );
buf1 gate1059( .a(N3453), .O(N3576) );
buf1 gate1060( .a(N3450), .O(N3579) );
buf1 gate1061( .a(N3459), .O(N3585) );
buf1 gate1062( .a(N3456), .O(N3588) );
inv1 gate1063( .a(N3522), .O(N3592) );
nand2 gate1064( .a(N3522), .b(N3405), .O(N3593) );
inv1 gate1065( .a(N3525), .O(N3594) );
nand2 gate1066( .a(N3525), .b(N3406), .O(N3595) );
inv1 gate1067( .a(N3528), .O(N3596) );
inv1 gate( .a(N3528),.O(N3528_NOT) );
inv1 gate( .a(N2630),.O(N2630_NOT));
and2 gate( .a(N3528_NOT), .b(p329), .O(EX821) );
and2 gate( .a(N2630_NOT), .b(EX821), .O(EX822) );
and2 gate( .a(N3528), .b(p330), .O(EX823) );
and2 gate( .a(N2630_NOT), .b(EX823), .O(EX824) );
and2 gate( .a(N3528_NOT), .b(p331), .O(EX825) );
and2 gate( .a(N2630), .b(EX825), .O(EX826) );
and2 gate( .a(N3528), .b(p332), .O(EX827) );
and2 gate( .a(N2630), .b(EX827), .O(EX828) );
or2  gate( .a(EX822), .b(EX824), .O(EX829) );
or2  gate( .a(EX826), .b(EX829), .O(EX830) );
or2  gate( .a(EX828), .b(EX830), .O(N3597) );
inv1 gate( .a(N3531),.O(N3531_NOT) );
inv1 gate( .a(N2376),.O(N2376_NOT));
and2 gate( .a(N3531_NOT), .b(p333), .O(EX831) );
and2 gate( .a(N2376_NOT), .b(EX831), .O(EX832) );
and2 gate( .a(N3531), .b(p334), .O(EX833) );
and2 gate( .a(N2376_NOT), .b(EX833), .O(EX834) );
and2 gate( .a(N3531_NOT), .b(p335), .O(EX835) );
and2 gate( .a(N2376), .b(EX835), .O(EX836) );
and2 gate( .a(N3531), .b(p336), .O(EX837) );
and2 gate( .a(N2376), .b(EX837), .O(EX838) );
or2  gate( .a(EX832), .b(EX834), .O(EX839) );
or2  gate( .a(EX836), .b(EX839), .O(EX840) );
or2  gate( .a(EX838), .b(EX840), .O(N3598) );
inv1 gate1070( .a(N3531), .O(N3599) );
and2 gate1071( .a(N3551), .b(N800), .O(N3600) );
nand2 gate1072( .a(N3552), .b(N3483), .O(N3603) );
nand2 gate1073( .a(N3553), .b(N3485), .O(N3608) );
inv1 gate( .a(N3554),.O(N3554_NOT) );
inv1 gate( .a(N3487),.O(N3487_NOT));
and2 gate( .a(N3554_NOT), .b(p337), .O(EX841) );
and2 gate( .a(N3487_NOT), .b(EX841), .O(EX842) );
and2 gate( .a(N3554), .b(p338), .O(EX843) );
and2 gate( .a(N3487_NOT), .b(EX843), .O(EX844) );
and2 gate( .a(N3554_NOT), .b(p339), .O(EX845) );
and2 gate( .a(N3487), .b(EX845), .O(EX846) );
and2 gate( .a(N3554), .b(p340), .O(EX847) );
and2 gate( .a(N3487), .b(EX847), .O(EX848) );
or2  gate( .a(EX842), .b(EX844), .O(EX849) );
or2  gate( .a(EX846), .b(EX849), .O(EX850) );
or2  gate( .a(EX848), .b(EX850), .O(N3612) );
inv1 gate( .a(N3555),.O(N3555_NOT) );
inv1 gate( .a(N3489),.O(N3489_NOT));
and2 gate( .a(N3555_NOT), .b(p341), .O(EX851) );
and2 gate( .a(N3489_NOT), .b(EX851), .O(EX852) );
and2 gate( .a(N3555), .b(p342), .O(EX853) );
and2 gate( .a(N3489_NOT), .b(EX853), .O(EX854) );
and2 gate( .a(N3555_NOT), .b(p343), .O(EX855) );
and2 gate( .a(N3489), .b(EX855), .O(EX856) );
and2 gate( .a(N3555), .b(p344), .O(EX857) );
and2 gate( .a(N3489), .b(EX857), .O(EX858) );
or2  gate( .a(EX852), .b(EX854), .O(EX859) );
or2  gate( .a(EX856), .b(EX859), .O(EX860) );
or2  gate( .a(EX858), .b(EX860), .O(N3615) );
inv1 gate( .a(N3556),.O(N3556_NOT) );
inv1 gate( .a(N3491),.O(N3491_NOT));
and2 gate( .a(N3556_NOT), .b(p345), .O(EX861) );
and2 gate( .a(N3491_NOT), .b(EX861), .O(EX862) );
and2 gate( .a(N3556), .b(p346), .O(EX863) );
and2 gate( .a(N3491_NOT), .b(EX863), .O(EX864) );
and2 gate( .a(N3556_NOT), .b(p347), .O(EX865) );
and2 gate( .a(N3491), .b(EX865), .O(EX866) );
and2 gate( .a(N3556), .b(p348), .O(EX867) );
and2 gate( .a(N3491), .b(EX867), .O(EX868) );
or2  gate( .a(EX862), .b(EX864), .O(EX869) );
or2  gate( .a(EX866), .b(EX869), .O(EX870) );
or2  gate( .a(EX868), .b(EX870), .O(N3616) );
nand2 gate1077( .a(N3557), .b(N3493), .O(N3622) );
inv1 gate1078( .a(N3534), .O(N3629) );
nand2 gate1079( .a(N3534), .b(N2645), .O(N3630) );
inv1 gate1080( .a(N3537), .O(N3631) );
inv1 gate( .a(N3537),.O(N3537_NOT) );
inv1 gate( .a(N2655),.O(N2655_NOT));
and2 gate( .a(N3537_NOT), .b(p349), .O(EX871) );
and2 gate( .a(N2655_NOT), .b(EX871), .O(EX872) );
and2 gate( .a(N3537), .b(p350), .O(EX873) );
and2 gate( .a(N2655_NOT), .b(EX873), .O(EX874) );
and2 gate( .a(N3537_NOT), .b(p351), .O(EX875) );
and2 gate( .a(N2655), .b(EX875), .O(EX876) );
and2 gate( .a(N3537), .b(p352), .O(EX877) );
and2 gate( .a(N2655), .b(EX877), .O(EX878) );
or2  gate( .a(EX872), .b(EX874), .O(EX879) );
or2  gate( .a(EX876), .b(EX879), .O(EX880) );
or2  gate( .a(EX878), .b(EX880), .O(N3632) );
nand2 gate1082( .a(N3540), .b(N2403), .O(N3633) );
inv1 gate1083( .a(N3540), .O(N3634) );
nand2 gate1084( .a(N3563), .b(N3502), .O(N3635) );
inv1 gate( .a(N3564),.O(N3564_NOT) );
inv1 gate( .a(N3504),.O(N3504_NOT));
and2 gate( .a(N3564_NOT), .b(p353), .O(EX881) );
and2 gate( .a(N3504_NOT), .b(EX881), .O(EX882) );
and2 gate( .a(N3564), .b(p354), .O(EX883) );
and2 gate( .a(N3504_NOT), .b(EX883), .O(EX884) );
and2 gate( .a(N3564_NOT), .b(p355), .O(EX885) );
and2 gate( .a(N3504), .b(EX885), .O(EX886) );
and2 gate( .a(N3564), .b(p356), .O(EX887) );
and2 gate( .a(N3504), .b(EX887), .O(EX888) );
or2  gate( .a(EX882), .b(EX884), .O(EX889) );
or2  gate( .a(EX886), .b(EX889), .O(EX890) );
or2  gate( .a(EX888), .b(EX890), .O(N3640) );
nand2 gate1086( .a(N3565), .b(N3506), .O(N3644) );
nand2 gate1087( .a(N3566), .b(N3508), .O(N3647) );
nand2 gate1088( .a(N3567), .b(N3510), .O(N3648) );
nand2 gate1089( .a(N3568), .b(N3512), .O(N3654) );
inv1 gate1090( .a(N3543), .O(N3661) );
nand2 gate1091( .a(N3543), .b(N2656), .O(N3662) );
inv1 gate( .a(N3238),.O(N3238_NOT) );
inv1 gate( .a(N3592),.O(N3592_NOT));
and2 gate( .a(N3238_NOT), .b(p357), .O(EX891) );
and2 gate( .a(N3592_NOT), .b(EX891), .O(EX892) );
and2 gate( .a(N3238), .b(p358), .O(EX893) );
and2 gate( .a(N3592_NOT), .b(EX893), .O(EX894) );
and2 gate( .a(N3238_NOT), .b(p359), .O(EX895) );
and2 gate( .a(N3592), .b(EX895), .O(EX896) );
and2 gate( .a(N3238), .b(p360), .O(EX897) );
and2 gate( .a(N3592), .b(EX897), .O(EX898) );
or2  gate( .a(EX892), .b(EX894), .O(EX899) );
or2  gate( .a(EX896), .b(EX899), .O(EX900) );
or2  gate( .a(EX898), .b(EX900), .O(N3667) );
nand2 gate1093( .a(N3241), .b(N3594), .O(N3668) );
nand2 gate1094( .a(N2472), .b(N3596), .O(N3669) );
nand2 gate1095( .a(N2213), .b(N3599), .O(N3670) );
buf1 gate1096( .a(N3600), .O(N3671) );
inv1 gate1097( .a(N3576), .O(N3691) );
inv1 gate( .a(N3576),.O(N3576_NOT) );
inv1 gate( .a(N3494),.O(N3494_NOT));
and2 gate( .a(N3576_NOT), .b(p361), .O(EX901) );
and2 gate( .a(N3494_NOT), .b(EX901), .O(EX902) );
and2 gate( .a(N3576), .b(p362), .O(EX903) );
and2 gate( .a(N3494_NOT), .b(EX903), .O(EX904) );
and2 gate( .a(N3576_NOT), .b(p363), .O(EX905) );
and2 gate( .a(N3494), .b(EX905), .O(EX906) );
and2 gate( .a(N3576), .b(p364), .O(EX907) );
and2 gate( .a(N3494), .b(EX907), .O(EX908) );
or2  gate( .a(EX902), .b(EX904), .O(EX909) );
or2  gate( .a(EX906), .b(EX909), .O(EX910) );
or2  gate( .a(EX908), .b(EX910), .O(N3692) );
inv1 gate1099( .a(N3579), .O(N3693) );
nand2 gate1100( .a(N3579), .b(N3496), .O(N3694) );
nand2 gate1101( .a(N2475), .b(N3629), .O(N3695) );
nand2 gate1102( .a(N2478), .b(N3631), .O(N3696) );
nand2 gate1103( .a(N2216), .b(N3634), .O(N3697) );
inv1 gate1104( .a(N3585), .O(N3716) );
nand2 gate1105( .a(N3585), .b(N3513), .O(N3717) );
inv1 gate1106( .a(N3588), .O(N3718) );
nand2 gate1107( .a(N3588), .b(N3515), .O(N3719) );
nand2 gate1108( .a(N2481), .b(N3661), .O(N3720) );
nand2 gate1109( .a(N3667), .b(N3593), .O(N3721) );
nand2 gate1110( .a(N3668), .b(N3595), .O(N3722) );
nand2 gate1111( .a(N3669), .b(N3597), .O(N3723) );
nand2 gate1112( .a(N3670), .b(N3598), .O(N3726) );
inv1 gate1113( .a(N3600), .O(N3727) );
nand2 gate1114( .a(N3364), .b(N3691), .O(N3728) );
nand2 gate1115( .a(N3367), .b(N3693), .O(N3729) );
nand2 gate1116( .a(N3695), .b(N3630), .O(N3730) );
and4 gate1117( .a(N3608), .b(N3615), .c(N3612), .d(N3603), .O(N3731) );
and2 gate1118( .a(N3603), .b(N3293), .O(N3732) );
and3 gate1119( .a(N3608), .b(N3603), .c(N3295), .O(N3733) );
and4 gate1120( .a(N3612), .b(N3603), .c(N3296), .d(N3608), .O(N3734) );
and2 gate1121( .a(N3616), .b(N3301), .O(N3735) );
and3 gate1122( .a(N3622), .b(N3616), .c(N3558), .O(N3736) );
nand2 gate1123( .a(N3696), .b(N3632), .O(N3737) );
nand2 gate1124( .a(N3697), .b(N3633), .O(N3740) );
nand2 gate1125( .a(N3394), .b(N3716), .O(N3741) );
nand2 gate1126( .a(N3397), .b(N3718), .O(N3742) );
nand2 gate1127( .a(N3720), .b(N3662), .O(N3743) );
and4 gate1128( .a(N3640), .b(N3647), .c(N3644), .d(N3635), .O(N3744) );
and2 gate1129( .a(N3635), .b(N3306), .O(N3745) );
and3 gate1130( .a(N3640), .b(N3635), .c(N3308), .O(N3746) );
and4 gate1131( .a(N3644), .b(N3635), .c(N3309), .d(N3640), .O(N3747) );
and2 gate1132( .a(N3648), .b(N3314), .O(N3748) );
and3 gate1133( .a(N3654), .b(N3648), .c(N3569), .O(N3749) );
inv1 gate1134( .a(N3721), .O(N3750) );
and2 gate1135( .a(N3722), .b(N246), .O(N3753) );
nand2 gate1136( .a(N3728), .b(N3692), .O(N3754) );
inv1 gate( .a(N3729),.O(N3729_NOT) );
inv1 gate( .a(N3694),.O(N3694_NOT));
and2 gate( .a(N3729_NOT), .b(p365), .O(EX911) );
and2 gate( .a(N3694_NOT), .b(EX911), .O(EX912) );
and2 gate( .a(N3729), .b(p366), .O(EX913) );
and2 gate( .a(N3694_NOT), .b(EX913), .O(EX914) );
and2 gate( .a(N3729_NOT), .b(p367), .O(EX915) );
and2 gate( .a(N3694), .b(EX915), .O(EX916) );
and2 gate( .a(N3729), .b(p368), .O(EX917) );
and2 gate( .a(N3694), .b(EX917), .O(EX918) );
or2  gate( .a(EX912), .b(EX914), .O(EX919) );
or2  gate( .a(EX916), .b(EX919), .O(EX920) );
or2  gate( .a(EX918), .b(EX920), .O(N3758) );
inv1 gate1138( .a(N3731), .O(N3761) );
or4 gate1139( .a(N3291), .b(N3732), .c(N3733), .d(N3734), .O(N3762) );
nand2 gate1140( .a(N3741), .b(N3717), .O(N3767) );
nand2 gate1141( .a(N3742), .b(N3719), .O(N3771) );
inv1 gate1142( .a(N3744), .O(N3774) );
or4 gate1143( .a(N3304), .b(N3745), .c(N3746), .d(N3747), .O(N3775) );
and2 gate1144( .a(N3723), .b(N3480), .O(N3778) );
and3 gate1145( .a(N3726), .b(N3723), .c(N3409), .O(N3779) );
or2 gate1146( .a(N2125), .b(N3753), .O(N3780) );
and2 gate1147( .a(N3750), .b(N800), .O(N3790) );
inv1 gate( .a(N3737),.O(N3737_NOT) );
inv1 gate( .a(N3500),.O(N3500_NOT));
and2 gate( .a(N3737_NOT), .b(p369), .O(EX921) );
and2 gate( .a(N3500_NOT), .b(EX921), .O(EX922) );
and2 gate( .a(N3737), .b(p370), .O(EX923) );
and2 gate( .a(N3500_NOT), .b(EX923), .O(EX924) );
and2 gate( .a(N3737_NOT), .b(p371), .O(EX925) );
and2 gate( .a(N3500), .b(EX925), .O(EX926) );
and2 gate( .a(N3737), .b(p372), .O(EX927) );
and2 gate( .a(N3500), .b(EX927), .O(EX928) );
or2  gate( .a(EX922), .b(EX924), .O(EX929) );
or2  gate( .a(EX926), .b(EX929), .O(EX930) );
or2  gate( .a(EX928), .b(EX930), .O(N3793) );
and3 gate1149( .a(N3740), .b(N3737), .c(N3428), .O(N3794) );
or3 gate1150( .a(N3479), .b(N3778), .c(N3779), .O(N3802) );
buf1 gate1151( .a(N3780), .O(N3803) );
buf1 gate1152( .a(N3780), .O(N3804) );
inv1 gate1153( .a(N3762), .O(N3805) );
and5 gate1154( .a(N3622), .b(N3730), .c(N3754), .d(N3616), .e(N3758), .O(N3806) );
and4 gate1155( .a(N3754), .b(N3616), .c(N3559), .d(N3622), .O(N3807) );
and5 gate1156( .a(N3758), .b(N3754), .c(N3616), .d(N3498), .e(N3622), .O(N3808) );
buf1 gate1157( .a(N3790), .O(N3809) );
or3 gate1158( .a(N3499), .b(N3793), .c(N3794), .O(N3811) );
inv1 gate1159( .a(N3775), .O(N3812) );
and5 gate1160( .a(N3654), .b(N3743), .c(N3767), .d(N3648), .e(N3771), .O(N3813) );
and4 gate1161( .a(N3767), .b(N3648), .c(N3570), .d(N3654), .O(N3814) );
and5 gate1162( .a(N3771), .b(N3767), .c(N3648), .d(N3517), .e(N3654), .O(N3815) );
or5 gate1163( .a(N3299), .b(N3735), .c(N3736), .d(N3807), .e(N3808), .O(N3816) );
and2 gate1164( .a(N3806), .b(N3802), .O(N3817) );
nand2 gate1165( .a(N3805), .b(N3761), .O(N3818) );
inv1 gate1166( .a(N3790), .O(N3819) );
or5 gate1167( .a(N3312), .b(N3748), .c(N3749), .d(N3814), .e(N3815), .O(N3820) );
and2 gate1168( .a(N3813), .b(N3811), .O(N3821) );
nand2 gate1169( .a(N3812), .b(N3774), .O(N3822) );
inv1 gate( .a(N3816),.O(N3816_NOT) );
inv1 gate( .a(N3817),.O(N3817_NOT));
and2 gate( .a(N3816_NOT), .b(p373), .O(EX931) );
and2 gate( .a(N3817_NOT), .b(EX931), .O(EX932) );
and2 gate( .a(N3816), .b(p374), .O(EX933) );
and2 gate( .a(N3817_NOT), .b(EX933), .O(EX934) );
and2 gate( .a(N3816_NOT), .b(p375), .O(EX935) );
and2 gate( .a(N3817), .b(EX935), .O(EX936) );
and2 gate( .a(N3816), .b(p376), .O(EX937) );
and2 gate( .a(N3817), .b(EX937), .O(EX938) );
or2  gate( .a(EX932), .b(EX934), .O(EX939) );
or2  gate( .a(EX936), .b(EX939), .O(EX940) );
or2  gate( .a(EX938), .b(EX940), .O(N3823) );
and3 gate1171( .a(N3727), .b(N3819), .c(N2841), .O(N3826) );
or2 gate1172( .a(N3820), .b(N3821), .O(N3827) );
inv1 gate1173( .a(N3823), .O(N3834) );
inv1 gate( .a(N3818),.O(N3818_NOT) );
inv1 gate( .a(N3823),.O(N3823_NOT));
and2 gate( .a(N3818_NOT), .b(p377), .O(EX941) );
and2 gate( .a(N3823_NOT), .b(EX941), .O(EX942) );
and2 gate( .a(N3818), .b(p378), .O(EX943) );
and2 gate( .a(N3823_NOT), .b(EX943), .O(EX944) );
and2 gate( .a(N3818_NOT), .b(p379), .O(EX945) );
and2 gate( .a(N3823), .b(EX945), .O(EX946) );
and2 gate( .a(N3818), .b(p380), .O(EX947) );
and2 gate( .a(N3823), .b(EX947), .O(EX948) );
or2  gate( .a(EX942), .b(EX944), .O(EX949) );
or2  gate( .a(EX946), .b(EX949), .O(EX950) );
or2  gate( .a(EX948), .b(EX950), .O(N3835) );
inv1 gate1175( .a(N3827), .O(N3836) );
and2 gate1176( .a(N3822), .b(N3827), .O(N3837) );
and2 gate1177( .a(N3762), .b(N3834), .O(N3838) );
and2 gate1178( .a(N3775), .b(N3836), .O(N3839) );
or2 gate1179( .a(N3838), .b(N3835), .O(N3840) );
or2 gate1180( .a(N3839), .b(N3837), .O(N3843) );
buf1 gate1181( .a(N3843), .O(N3851) );
nand2 gate1182( .a(N3843), .b(N3840), .O(N3852) );
and2 gate1183( .a(N3843), .b(N3852), .O(N3857) );
and2 gate1184( .a(N3852), .b(N3840), .O(N3858) );
or2 gate1185( .a(N3857), .b(N3858), .O(N3859) );
inv1 gate1186( .a(N3859), .O(N3864) );
and2 gate1187( .a(N3859), .b(N3864), .O(N3869) );
or2 gate1188( .a(N3869), .b(N3864), .O(N3870) );
inv1 gate1189( .a(N3870), .O(N3875) );
and3 gate1190( .a(N2826), .b(N3028), .c(N3870), .O(N3876) );
and3 gate1191( .a(N3826), .b(N3876), .c(N1591), .O(N3877) );
buf1 gate1192( .a(N3877), .O(N3881) );
inv1 gate1193( .a(N3877), .O(N3882) );
buf1 gate1194( .a(N143_I), .O(N143_O) );
buf1 gate1195( .a(N144_I), .O(N144_O) );
buf1 gate1196( .a(N145_I), .O(N145_O) );
buf1 gate1197( .a(N146_I), .O(N146_O) );
buf1 gate1198( .a(N147_I), .O(N147_O) );
buf1 gate1199( .a(N148_I), .O(N148_O) );
buf1 gate1200( .a(N149_I), .O(N149_O) );
buf1 gate1201( .a(N150_I), .O(N150_O) );
buf1 gate1202( .a(N151_I), .O(N151_O) );
buf1 gate1203( .a(N152_I), .O(N152_O) );
buf1 gate1204( .a(N153_I), .O(N153_O) );
buf1 gate1205( .a(N154_I), .O(N154_O) );
buf1 gate1206( .a(N155_I), .O(N155_O) );
buf1 gate1207( .a(N156_I), .O(N156_O) );
buf1 gate1208( .a(N157_I), .O(N157_O) );
buf1 gate1209( .a(N158_I), .O(N158_O) );
buf1 gate1210( .a(N159_I), .O(N159_O) );
buf1 gate1211( .a(N160_I), .O(N160_O) );
buf1 gate1212( .a(N161_I), .O(N161_O) );
buf1 gate1213( .a(N162_I), .O(N162_O) );
buf1 gate1214( .a(N163_I), .O(N163_O) );
buf1 gate1215( .a(N164_I), .O(N164_O) );
buf1 gate1216( .a(N165_I), .O(N165_O) );
buf1 gate1217( .a(N166_I), .O(N166_O) );
buf1 gate1218( .a(N167_I), .O(N167_O) );
buf1 gate1219( .a(N168_I), .O(N168_O) );
buf1 gate1220( .a(N169_I), .O(N169_O) );
buf1 gate1221( .a(N170_I), .O(N170_O) );
buf1 gate1222( .a(N171_I), .O(N171_O) );
buf1 gate1223( .a(N172_I), .O(N172_O) );
buf1 gate1224( .a(N173_I), .O(N173_O) );
buf1 gate1225( .a(N174_I), .O(N174_O) );
buf1 gate1226( .a(N175_I), .O(N175_O) );
buf1 gate1227( .a(N176_I), .O(N176_O) );
buf1 gate1228( .a(N177_I), .O(N177_O) );
buf1 gate1229( .a(N178_I), .O(N178_O) );
buf1 gate1230( .a(N179_I), .O(N179_O) );
buf1 gate1231( .a(N180_I), .O(N180_O) );
buf1 gate1232( .a(N181_I), .O(N181_O) );
buf1 gate1233( .a(N182_I), .O(N182_O) );
buf1 gate1234( .a(N183_I), .O(N183_O) );
buf1 gate1235( .a(N184_I), .O(N184_O) );
buf1 gate1236( .a(N185_I), .O(N185_O) );
buf1 gate1237( .a(N186_I), .O(N186_O) );
buf1 gate1238( .a(N187_I), .O(N187_O) );
buf1 gate1239( .a(N188_I), .O(N188_O) );
buf1 gate1240( .a(N189_I), .O(N189_O) );
buf1 gate1241( .a(N190_I), .O(N190_O) );
buf1 gate1242( .a(N191_I), .O(N191_O) );
buf1 gate1243( .a(N192_I), .O(N192_O) );
buf1 gate1244( .a(N193_I), .O(N193_O) );
buf1 gate1245( .a(N194_I), .O(N194_O) );
buf1 gate1246( .a(N195_I), .O(N195_O) );
buf1 gate1247( .a(N196_I), .O(N196_O) );
buf1 gate1248( .a(N197_I), .O(N197_O) );
buf1 gate1249( .a(N198_I), .O(N198_O) );
buf1 gate1250( .a(N199_I), .O(N199_O) );
buf1 gate1251( .a(N200_I), .O(N200_O) );
buf1 gate1252( .a(N201_I), .O(N201_O) );
buf1 gate1253( .a(N202_I), .O(N202_O) );
buf1 gate1254( .a(N203_I), .O(N203_O) );
buf1 gate1255( .a(N204_I), .O(N204_O) );
buf1 gate1256( .a(N205_I), .O(N205_O) );
buf1 gate1257( .a(N206_I), .O(N206_O) );
buf1 gate1258( .a(N207_I), .O(N207_O) );
buf1 gate1259( .a(N208_I), .O(N208_O) );
buf1 gate1260( .a(N209_I), .O(N209_O) );
buf1 gate1261( .a(N210_I), .O(N210_O) );
buf1 gate1262( .a(N211_I), .O(N211_O) );
buf1 gate1263( .a(N212_I), .O(N212_O) );
buf1 gate1264( .a(N213_I), .O(N213_O) );
buf1 gate1265( .a(N214_I), .O(N214_O) );
buf1 gate1266( .a(N215_I), .O(N215_O) );
buf1 gate1267( .a(N216_I), .O(N216_O) );
buf1 gate1268( .a(N217_I), .O(N217_O) );
buf1 gate1269( .a(N218_I), .O(N218_O) );

endmodule
