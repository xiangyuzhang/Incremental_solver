module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115; // anything
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41; //RE__ALLOW(00,01,10);
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12;


inv1 gate1( .a(N1), .O(N118) );  // anything
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );

  xor2  gate441(.a(N30), .b(N126), .O(gate23inter0));
  nand2 gate442(.a(gate23inter0), .b(s_40), .O(gate23inter1));
  and2  gate443(.a(N30), .b(N126), .O(gate23inter2));
  inv1  gate444(.a(s_40), .O(gate23inter3));
  inv1  gate445(.a(s_41), .O(gate23inter4));
  nand2 gate446(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate447(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate448(.a(N126), .O(gate23inter7));
  inv1  gate449(.a(N30), .O(gate23inter8));
  nand2 gate450(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate451(.a(s_41), .b(gate23inter3), .O(gate23inter10));
  nor2  gate452(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate453(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate454(.a(gate23inter12), .b(gate23inter1), .O(N162));
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );

  xor2  gate301(.a(N69), .b(N138), .O(gate26inter0));
  nand2 gate302(.a(gate26inter0), .b(s_20), .O(gate26inter1));
  and2  gate303(.a(N69), .b(N138), .O(gate26inter2));
  inv1  gate304(.a(s_20), .O(gate26inter3));
  inv1  gate305(.a(s_21), .O(gate26inter4));
  nand2 gate306(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate307(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate308(.a(N138), .O(gate26inter7));
  inv1  gate309(.a(N69), .O(gate26inter8));
  nand2 gate310(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate311(.a(s_21), .b(gate26inter3), .O(gate26inter10));
  nor2  gate312(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate313(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate314(.a(gate26inter12), .b(gate26inter1), .O(N171));

  xor2  gate399(.a(N82), .b(N142), .O(gate27inter0));
  nand2 gate400(.a(gate27inter0), .b(s_34), .O(gate27inter1));
  and2  gate401(.a(N82), .b(N142), .O(gate27inter2));
  inv1  gate402(.a(s_34), .O(gate27inter3));
  inv1  gate403(.a(s_35), .O(gate27inter4));
  nand2 gate404(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate405(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate406(.a(N142), .O(gate27inter7));
  inv1  gate407(.a(N82), .O(gate27inter8));
  nand2 gate408(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate409(.a(s_35), .b(gate27inter3), .O(gate27inter10));
  nor2  gate410(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate411(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate412(.a(gate27inter12), .b(gate27inter1), .O(N174));
nand2 gate28( .a(N146), .b(N95), .O(N177) );
nand2 gate29( .a(N150), .b(N108), .O(N180) );
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );

  xor2  gate287(.a(N131), .b(N47), .O(gate34inter0));
  nand2 gate288(.a(gate34inter0), .b(s_18), .O(gate34inter1));
  and2  gate289(.a(N131), .b(N47), .O(gate34inter2));
  inv1  gate290(.a(s_18), .O(gate34inter3));
  inv1  gate291(.a(s_19), .O(gate34inter4));
  nand2 gate292(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate293(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate294(.a(N47), .O(gate34inter7));
  inv1  gate295(.a(N131), .O(gate34inter8));
  nand2 gate296(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate297(.a(s_19), .b(gate34inter3), .O(gate34inter10));
  nor2  gate298(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate299(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate300(.a(gate34inter12), .b(gate34inter1), .O(N187));
nor2 gate35( .a(N53), .b(N131), .O(N188) );

  xor2  gate329(.a(N135), .b(N60), .O(gate36inter0));
  nand2 gate330(.a(gate36inter0), .b(s_24), .O(gate36inter1));
  and2  gate331(.a(N135), .b(N60), .O(gate36inter2));
  inv1  gate332(.a(s_24), .O(gate36inter3));
  inv1  gate333(.a(s_25), .O(gate36inter4));
  nand2 gate334(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate335(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate336(.a(N60), .O(gate36inter7));
  inv1  gate337(.a(N135), .O(gate36inter8));
  nand2 gate338(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate339(.a(s_25), .b(gate36inter3), .O(gate36inter10));
  nor2  gate340(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate341(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate342(.a(gate36inter12), .b(gate36inter1), .O(N189));
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );
nor2 gate41( .a(N92), .b(N143), .O(N194) );
nor2 gate42( .a(N99), .b(N147), .O(N195) );

  xor2  gate315(.a(N147), .b(N105), .O(gate43inter0));
  nand2 gate316(.a(gate43inter0), .b(s_22), .O(gate43inter1));
  and2  gate317(.a(N147), .b(N105), .O(gate43inter2));
  inv1  gate318(.a(s_22), .O(gate43inter3));
  inv1  gate319(.a(s_23), .O(gate43inter4));
  nand2 gate320(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate321(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate322(.a(N105), .O(gate43inter7));
  inv1  gate323(.a(N147), .O(gate43inter8));
  nand2 gate324(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate325(.a(s_23), .b(gate43inter3), .O(gate43inter10));
  nor2  gate326(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate327(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate328(.a(gate43inter12), .b(gate43inter1), .O(N196));
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );
xor2 gate52( .a(N203), .b(N162), .O(N230) );

  xor2  gate273(.a(N165), .b(N203), .O(gate53inter0));
  nand2 gate274(.a(gate53inter0), .b(s_16), .O(gate53inter1));
  and2  gate275(.a(N165), .b(N203), .O(gate53inter2));
  inv1  gate276(.a(s_16), .O(gate53inter3));
  inv1  gate277(.a(s_17), .O(gate53inter4));
  nand2 gate278(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate279(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate280(.a(N203), .O(gate53inter7));
  inv1  gate281(.a(N165), .O(gate53inter8));
  nand2 gate282(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate283(.a(s_17), .b(gate53inter3), .O(gate53inter10));
  nor2  gate284(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate285(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate286(.a(gate53inter12), .b(gate53inter1), .O(N233));

  xor2  gate175(.a(N168), .b(N203), .O(gate54inter0));
  nand2 gate176(.a(gate54inter0), .b(s_2), .O(gate54inter1));
  and2  gate177(.a(N168), .b(N203), .O(gate54inter2));
  inv1  gate178(.a(s_2), .O(gate54inter3));
  inv1  gate179(.a(s_3), .O(gate54inter4));
  nand2 gate180(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate181(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate182(.a(N203), .O(gate54inter7));
  inv1  gate183(.a(N168), .O(gate54inter8));
  nand2 gate184(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate185(.a(s_3), .b(gate54inter3), .O(gate54inter10));
  nor2  gate186(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate187(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate188(.a(gate54inter12), .b(gate54inter1), .O(N236));
xor2 gate55( .a(N203), .b(N171), .O(N239) );

  xor2  gate371(.a(N213), .b(N1), .O(gate56inter0));
  nand2 gate372(.a(gate56inter0), .b(s_30), .O(gate56inter1));
  and2  gate373(.a(N213), .b(N1), .O(gate56inter2));
  inv1  gate374(.a(s_30), .O(gate56inter3));
  inv1  gate375(.a(s_31), .O(gate56inter4));
  nand2 gate376(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate377(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate378(.a(N1), .O(gate56inter7));
  inv1  gate379(.a(N213), .O(gate56inter8));
  nand2 gate380(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate381(.a(s_31), .b(gate56inter3), .O(gate56inter10));
  nor2  gate382(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate383(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate384(.a(gate56inter12), .b(gate56inter1), .O(N242));
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );

  xor2  gate217(.a(N37), .b(N213), .O(gate62inter0));
  nand2 gate218(.a(gate62inter0), .b(s_8), .O(gate62inter1));
  and2  gate219(.a(N37), .b(N213), .O(gate62inter2));
  inv1  gate220(.a(s_8), .O(gate62inter3));
  inv1  gate221(.a(s_9), .O(gate62inter4));
  nand2 gate222(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate223(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate224(.a(N213), .O(gate62inter7));
  inv1  gate225(.a(N37), .O(gate62inter8));
  nand2 gate226(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate227(.a(s_9), .b(gate62inter3), .O(gate62inter10));
  nor2  gate228(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate229(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate230(.a(gate62inter12), .b(gate62inter1), .O(N254));
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );

  xor2  gate161(.a(N157), .b(N224), .O(gate68inter0));
  nand2 gate162(.a(gate68inter0), .b(s_0), .O(gate68inter1));
  and2  gate163(.a(N157), .b(N224), .O(gate68inter2));
  inv1  gate164(.a(s_0), .O(gate68inter3));
  inv1  gate165(.a(s_1), .O(gate68inter4));
  nand2 gate166(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate167(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate168(.a(N224), .O(gate68inter7));
  inv1  gate169(.a(N157), .O(gate68inter8));
  nand2 gate170(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate171(.a(s_1), .b(gate68inter3), .O(gate68inter10));
  nor2  gate172(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate173(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate174(.a(gate68inter12), .b(gate68inter1), .O(N260));
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );
nand2 gate71( .a(N230), .b(N185), .O(N267) );
nand2 gate72( .a(N233), .b(N187), .O(N270) );
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );

  xor2  gate385(.a(N184), .b(N227), .O(gate78inter0));
  nand2 gate386(.a(gate78inter0), .b(s_32), .O(gate78inter1));
  and2  gate387(.a(N184), .b(N227), .O(gate78inter2));
  inv1  gate388(.a(s_32), .O(gate78inter3));
  inv1  gate389(.a(s_33), .O(gate78inter4));
  nand2 gate390(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate391(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate392(.a(N227), .O(gate78inter7));
  inv1  gate393(.a(N184), .O(gate78inter8));
  nand2 gate394(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate395(.a(s_33), .b(gate78inter3), .O(gate78inter10));
  nor2  gate396(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate397(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate398(.a(gate78inter12), .b(gate78inter1), .O(N288));
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );

  xor2  gate231(.a(N194), .b(N243), .O(gate83inter0));
  nand2 gate232(.a(gate83inter0), .b(s_10), .O(gate83inter1));
  and2  gate233(.a(N194), .b(N243), .O(gate83inter2));
  inv1  gate234(.a(s_10), .O(gate83inter3));
  inv1  gate235(.a(s_11), .O(gate83inter4));
  nand2 gate236(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate237(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate238(.a(N243), .O(gate83inter7));
  inv1  gate239(.a(N194), .O(gate83inter8));
  nand2 gate240(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate241(.a(s_11), .b(gate83inter3), .O(gate83inter10));
  nor2  gate242(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate243(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate244(.a(gate83inter12), .b(gate83inter1), .O(N293));
nand2 gate84( .a(N247), .b(N196), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319), .b(N60), .O(N342) );

  xor2  gate203(.a(N285), .b(N309), .O(gate112inter0));
  nand2 gate204(.a(gate112inter0), .b(s_6), .O(gate112inter1));
  and2  gate205(.a(N285), .b(N309), .O(gate112inter2));
  inv1  gate206(.a(s_6), .O(gate112inter3));
  inv1  gate207(.a(s_7), .O(gate112inter4));
  nand2 gate208(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate209(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate210(.a(N309), .O(gate112inter7));
  inv1  gate211(.a(N285), .O(gate112inter8));
  nand2 gate212(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate213(.a(s_7), .b(gate112inter3), .O(gate112inter10));
  nor2  gate214(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate215(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate216(.a(gate112inter12), .b(gate112inter1), .O(N343));

  xor2  gate189(.a(N73), .b(N319), .O(gate113inter0));
  nand2 gate190(.a(gate113inter0), .b(s_4), .O(gate113inter1));
  and2  gate191(.a(N73), .b(N319), .O(gate113inter2));
  inv1  gate192(.a(s_4), .O(gate113inter3));
  inv1  gate193(.a(s_5), .O(gate113inter4));
  nand2 gate194(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate195(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate196(.a(N319), .O(gate113inter7));
  inv1  gate197(.a(N73), .O(gate113inter8));
  nand2 gate198(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate199(.a(s_5), .b(gate113inter3), .O(gate113inter10));
  nor2  gate200(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate201(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate202(.a(gate113inter12), .b(gate113inter1), .O(N344));

  xor2  gate343(.a(N86), .b(N319), .O(gate114inter0));
  nand2 gate344(.a(gate114inter0), .b(s_26), .O(gate114inter1));
  and2  gate345(.a(N86), .b(N319), .O(gate114inter2));
  inv1  gate346(.a(s_26), .O(gate114inter3));
  inv1  gate347(.a(s_27), .O(gate114inter4));
  nand2 gate348(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate349(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate350(.a(N319), .O(gate114inter7));
  inv1  gate351(.a(N86), .O(gate114inter8));
  nand2 gate352(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate353(.a(s_27), .b(gate114inter3), .O(gate114inter10));
  nor2  gate354(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate355(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate356(.a(gate114inter12), .b(gate114inter1), .O(N345));
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );

  xor2  gate357(.a(N300), .b(N330), .O(gate117inter0));
  nand2 gate358(.a(gate117inter0), .b(s_28), .O(gate117inter1));
  and2  gate359(.a(N300), .b(N330), .O(gate117inter2));
  inv1  gate360(.a(s_28), .O(gate117inter3));
  inv1  gate361(.a(s_29), .O(gate117inter4));
  nand2 gate362(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate363(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate364(.a(N330), .O(gate117inter7));
  inv1  gate365(.a(N300), .O(gate117inter8));
  nand2 gate366(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate367(.a(s_29), .b(gate117inter3), .O(gate117inter10));
  nor2  gate368(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate369(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate370(.a(gate117inter12), .b(gate117inter1), .O(N348));
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );

  xor2  gate413(.a(N303), .b(N333), .O(gate120inter0));
  nand2 gate414(.a(gate120inter0), .b(s_36), .O(gate120inter1));
  and2  gate415(.a(N303), .b(N333), .O(gate120inter2));
  inv1  gate416(.a(s_36), .O(gate120inter3));
  inv1  gate417(.a(s_37), .O(gate120inter4));
  nand2 gate418(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate419(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate420(.a(N333), .O(gate120inter7));
  inv1  gate421(.a(N303), .O(gate120inter8));
  nand2 gate422(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate423(.a(s_37), .b(gate120inter3), .O(gate120inter10));
  nor2  gate424(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate425(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate426(.a(gate120inter12), .b(gate120inter1), .O(N351));
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );

  xor2  gate259(.a(N27), .b(N360), .O(gate130inter0));
  nand2 gate260(.a(gate130inter0), .b(s_14), .O(gate130inter1));
  and2  gate261(.a(N27), .b(N360), .O(gate130inter2));
  inv1  gate262(.a(s_14), .O(gate130inter3));
  inv1  gate263(.a(s_15), .O(gate130inter4));
  nand2 gate264(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate265(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate266(.a(N360), .O(gate130inter7));
  inv1  gate267(.a(N27), .O(gate130inter8));
  nand2 gate268(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate269(.a(s_15), .b(gate130inter3), .O(gate130inter10));
  nor2  gate270(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate271(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate272(.a(gate130inter12), .b(gate130inter1), .O(N372));
nand2 gate131( .a(N360), .b(N40), .O(N373) );

  xor2  gate245(.a(N53), .b(N360), .O(gate132inter0));
  nand2 gate246(.a(gate132inter0), .b(s_12), .O(gate132inter1));
  and2  gate247(.a(N53), .b(N360), .O(gate132inter2));
  inv1  gate248(.a(s_12), .O(gate132inter3));
  inv1  gate249(.a(s_13), .O(gate132inter4));
  nand2 gate250(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate251(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate252(.a(N360), .O(gate132inter7));
  inv1  gate253(.a(N53), .O(gate132inter8));
  nand2 gate254(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate255(.a(s_13), .b(gate132inter3), .O(gate132inter10));
  nor2  gate256(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate257(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate258(.a(gate132inter12), .b(gate132inter1), .O(N374));
nand2 gate133( .a(N360), .b(N66), .O(N375) );

  xor2  gate427(.a(N79), .b(N360), .O(gate134inter0));
  nand2 gate428(.a(gate134inter0), .b(s_38), .O(gate134inter1));
  and2  gate429(.a(N79), .b(N360), .O(gate134inter2));
  inv1  gate430(.a(s_38), .O(gate134inter3));
  inv1  gate431(.a(s_39), .O(gate134inter4));
  nand2 gate432(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate433(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate434(.a(N360), .O(gate134inter7));
  inv1  gate435(.a(N79), .O(gate134inter8));
  nand2 gate436(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate437(.a(s_39), .b(gate134inter3), .O(gate134inter10));
  nor2  gate438(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate439(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate440(.a(gate134inter12), .b(gate134inter1), .O(N376));
nand2 gate135( .a(N360), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule
